// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
LoufMElIzLEs9F+po1uJxjBPw0zjiWmhh/xA3P+J0i807XjCbk8DQcBcoo8w0YvN
cNoEQoYuOolSIcuFlIlQIUzdFRxEEZEr/BzDUUCjZlUTY334iVcJZMj4yHRwmKSb
DdjZRypTHte6/acRzlFsO8BD22YFNaMBZ691Lvh14OqLT0gQ4+9Trw==
//pragma protect end_key_block
//pragma protect digest_block
UJtf9bqIoZa28Fzhqh8tF1XubMw=
//pragma protect end_digest_block
//pragma protect data_block
BREprGEIEEIoksSsTjwuMCSVXqT+MyhEyBXebVb1SIpC7CIrzLwrtBIwCLRigPb+
XBfAcA2G4i0BZQUJMvK+rcBDqB0T3tUK/DiNgjufR2eBw1iGZEa5MwYUWYP1bKqM
/+Xe8B+Q7FPjJthU46w6iuoKFenEjebobRX9m47qACHk1jZnS6rYiXfjo9l3l536
Ifn5dsucseEP+tv2uDydUEZiQ0672MVTmOX9x2jSy3DXUUPmuelaOihqayv0SMdR
D4Xl8+6YUNIpLBcK6D1rn6U3Ql3uUJ+bCnV5S8ACcz3rhVuLXp/BIVFo0DfeXqJJ
2ikYC5uaECWArrdhbVffK/f8lerTqVM69MrAMb20Mg8D6vN6fX4hNxNsa7a8ucaK
hzVXZ6CiEyG2PWirs5/gVfk/MbCfw6uITMUCegxRVm3CyibmFNF2BTe55e4WQkru
fZi/AvxD9g5/fzzADXL6b/PvdtCq2afPRyjsufK6/EvoQ96w7pPYHaXCkaklwkB6
F6VIY/benAIaqEVVjodJJv7gVJJ5zulqj1dIJzPlUmzeo6Nc67MeDa7OD7cOi804
earoyviQka6LLnCELJmsZ29s8ICqmxwrDoj3W1J6mz89oLJflnlfB5RIAo6ak19D
enFzZrejm1HoM4qgHEfhAECCV18z4V2w3sfpy1KDp/zBdBDxJ6e2mka6hEpO8fC+
7eZ530GVsaD0ILiXb5/NKleDdKzAu3xVc9ecQuQx3jbhQsMijrfD9moAqqrzYCN6
J8J4NYXC5YkcqILVhmsTOeAJ9vwD7GPftpnndYSowizq6UlXbK4ejLylUyDWClvU
GkDxRsSvvNh3LR5MBTX9lbsnkZO3NOnA9zCSywomYM+NtnTUyLAvijS95PuiWPNA
iuqMhGlMhlAvzFzzcR6B66/9iIK5XF8rFTIMLZt2YvC6yqnhRL7TU7t7ikVAyqvW
go9Br0stc9Mfcq07U3NslWDt0K/dpBzDo0FqgkNF2g3B2mYCdttIiZldAu/QuMSZ
nwKIWN6eQi0S+n3EJRxfdrKRintVJeUCwTJyhhtZU7ijVXwrQCiCZD6yRrFhlx0M
WHTcud4AVEWmvczQnlDPRZ3mUoJjzpzbKUrT88lsKpvi2olXg47A5i1o8a4RHu43
XXM1DPs2nJIdG5SWKHH0Wmg4UDmcmQNygpACZLLxxm9J/dYy/GRx/MHbN+n6/FZQ
SDvHmHZsiiwhDurjJvZIVHCXvsPfiVRVR++u/SXgUceE26c2TCDaasFsmCjRQMgA
rXvuxL6MRgshg6dl1UhW73LMMsxPHAzysWIDPGLsrOcdFBiGA/iaDJqJVNlzMclz
p9MTrSRHJkVwQXXk8eAu35KLi2G4xZQxagqD8TjG2yr8dsGnXU44ug6MXvm1Vj+M
qApBJzahhctt+YuE3+J1ae7TTv7139cBBBUfMLp/o/3yMBFV11zXUAKHztriVuNc
wW/eTIju+c0PD1yAMunfb1FJ2V+7qmyvdgF8oYLqDSq+WKaMgOIWuTjO2a1r9f5R
E5rJBq/rzHalcaDPFWjx0s7e5gwkRDr5XSyuRYA9/S4ugEgbCJcke+MF2uvcJk95
RemSsKdz1Aw1Rg3Q20bpK7W0JGsX+dw2QG0vKMkgDIzJx7SaTFTy6HZ3wyPxqWY3
cMI5vDnkO2gZMwQvKjdmZZLT8rdDKtpcrLZFIBrXT1b0nDES40FSo8xSGNQjB0k5
9vSya+SLnG4vjEWCyFvcag+IZycDEJrZcOHjsUyo988jOg3CjYYVaZvav65UoFur
Yr8IcP4XBrr6V2QmqnRUKS/sBNlg3TvUacJGhJRYZpAbgVUs2oeh16XNWoMtlqqA
SEVirFjZnhNgEAoddc4m6Tg3iavEz+qvSo3M+wv98AjbWIzKiuqxmNd6t9klq/iR
j7UE1bkYrXd2SWHWn4zwRUk45eYfryb6M2+sjpp6clPETo/zCTng4sTH5UqIeREH
c+ab9tb+HtH8vY9KuvvEnbq4obFe78nLQUCKQSmDrNO2VrqJstaKKrcDpHCNiuhx
XL/qhzy7iL5FGgqZPivp6dvNTQDvVhBvSqYqyvI+iUMPndD9/mlCLRx+yCTFMF0k
/sikvJyPy8uMrlnfBRILZZI/bBJi60G3kOy8vDeJgFrQ7YtS1k12j7m0lF/b/49S
5G4aKgxkeDJO9yxmrR6by+VGY7YTFs7YGRYzYPAG2kfyUgBzyi6WdWYyoKWKgksT
Wq0xu390IPVCPSgFzWJJjsmTAJaNGBl+0HtIJI7+X+J5plAfS8zBhJdupn3Jh6yp
iX1bSHH+PDJnPW6cMd28KJcQJKeE10XSQuRUcSkNe4b4zgAHyvGbf9PSLpEaBUpt
rxFg8OjPbsTiulZtoLK1HrMzm2U0Bj1ZBsivWrkftxhyEQLXM1/1ne5AzzL6eOi9
0g/5pO6y2KZPU+JBObA+Q8JGYcd1o+QdjHRfvp5EqCXSkLDt8vnOfplUuDdtCQZ/
hgKXdBxtGltEn3GuYpQLla5mOxingk0WBkCsipbhShw8avKnwrX5R2En7TruD0WW
67epTJH+wlIJ4OAy+o4RFjEHOuZLvkOj4vdmNAhiwTyDKuSAL5/OnbtH7z6oDqfo
QWDLkdKRD5ynifG6CN2wnLEcD4E7IAO1+r7JcfODRD+m6rTuYhpgMPehudQxcY/T
sb6FQ1O4IPoRDxLbqWpUTyz+PFFBBgxmXYdo3RVdWluP8BKIbhOBhPCmnORNuiZq
QZAll8vSaGG2Km0TQk/cXhfFm8emv9TibDAg2axpynB9JSEJ9QQ7UUmtvXLek9Ei
xbVyYcAy8yCGf5bHp/SxZJ2OONrEqEnJ6YuHP5Iwbt75sPkF2e/UY9I8MjMpKGPC
EZ5kAYtH20EuYmyTT/EkAkmRHc+jZlKf4prWupjYSFyjPCu1Pdv1/iAIyC5mKn++
vs6nesLfnPnNwAGi38JLzwDVb+3mMyHVj53iPqzSj9V0dBUHadxYY7pEWc04c4bw
zfxaNaNglkiL6vziDAi2jHtNUaqS0VcmpdQxLctCSwSg/sytVDhlkTv8y08cgTn1
FeOco43kV57LE0AN0HGFZHUJITL/8IdOd9pcUmoycUuGgndhKdhpjOsbFDAf615J
Mqej20pKggjdOHxRfZH4YA6brz8nqe1SxMfuGbV4+qi0OQ4fMpnMFivCScSTG54i
B3sqL0zHzUm+PN702UstubOTQZhVuogDu1o6/+srD5wNVYutCLAxo1JJf2OGZdct
0Pz+mGJjXniQB2mXo7HraMCDuNL2JGxlQH3o9F5bl2yc42WBz+nMxSlrItiFoi3u
oA2nAY218P/HXD5mXS0+hZ5x1JLb67lR/AtLHtUQNuOkjI3U1+LrUeUFiuijVyeZ
K5NYyhNPmtwJqdgWrsxOdtSDgi0y66dr8El8SN3AY5IeCed+cZ9k4+ldgl8+BeDw
nLw39BiMX7imWiOpKhAiflBjHwkUxe4Yp5GJXJoF5eR+KUe2yzYBtneO2thE9OAz
1AOtrm++/cyVFlPGluDnnS79sTKX7m11oIO6LC+t7YfnqY60fJyVRHmG93JnTWwz
BTeBfaf0yE34mWtU6XqjUQ0+2Zrpu8bzqb4EsRqwSS0QrjCS8tWLE6q0kfm5C3Kk
SxrN+OCopOrZ55sVJuz2DpwselbhFBQ00MEFvIg+7DAmZDnLm7WTrWz6q6q22I/s
X2KSB9HrYKynYPcFMbi/RkbRmmZnJ8Mmt+L+iJMrmqE+z3NJxknqtX8czE4/EDL/
d4iYd8nSLlNX/jWk6PHK4zoQk19f1MLbN22h7Y2CqFOno8JRp/Le2ucUg2b/fg2N
k7Kttu8W/rPu+gkaEzTjLDcEUx0WW90P+veERzSK5BV3dvNgkSQAPO65fkElfZdh
aDC927TuOUPjmGPMKCDEYgleO/eGDdqTnTW7N5qPcBT2SNFg5f2OhkoC6qfVsOje
e8U+uF04SBTFFFbocGD392l59xVdR4SKG7VW7YxtNF4dNsQGkNKl5GHjEW7zudBF
ImL9AoZ/is13LHGGer6w9VXb9JB+aICCjSTWF0iPs2pUwFJBR+M/a/6TeIxY2C7f
1lpWWr7IrMT7G92IviOMo8KDwuUqYEkf2k8VGUMbQFDnzs8TPdSRppZn9PfY6nL0
j9XeKxaaevZeuo6DXaijkh/WaiZfzNOlMjVbgVGVUtprjDeZM4AvrLKfJWsndddy
njgBP62MninoY6U2q0qrVpzTYNCoE8BYVFjksaLeqVHtMn4zDhUcc8w3FlzGEXXt
iSxd66wnH7aHAK4JNfWCv17yJYrXOJlTi5SBDv0tIhkJ6/kmtnGRs1uDLEH0u4vW
+UHzGhI35qz8CkvpL28JUZjg+hVbulrJJuQqB0dNeLes8PDBIyXxYEPXcx7n3VBk
OVbPrDrmcJvjMr89L1Cg6tYTR7a+ZU4MO0psfASvjQw5MMBB6Y6V0NfoSykilAiE
Nf2/cQZOYVDOVBWycTmJpP0JH4chCK7lNPUsEEgdafE931CUm/HbtMwTH9SfD0MW
GDoRRJ4ZRmfL4btrIuEBWSbMFU7jubtAIq8k7Ov9uAECZZoqhrrXhuFmLS+25GBS
EI2RLSvt6Og/OLAiJcHWtqa3tA1td4CW2yWPHrdRmfTVzTKZgWtu+r30aK0RgvNf
+wnQKrpXx4jqbHIambt+wLPEhH3BbwLGm4xI+42xRXJVc/7F1PN/mvgszsFSNFHP
O78erZe3PGhflS/VYeLHyHWdY2uim/x+Xk986pHhdV2M2CdM3nYBFXmwp+QG4FSc
J8RB/Gja/J+xVnNT5BCYg2hYZU7TXj+qBJqjObe/ARVw+YscHY3p9g28mE/AIxjh
qHdKz+0JAd5ENygd8m1wPlJvcIn/e/ngzFs5E48yB9021NWIkAS1V0pU/JHjX6J/
4E6Muhm0M2W3Cyhq5OADO4sml+fRrVcIPZ2/6K1vJWP9/O1OvT982OARGWsuMAyR
q1dSsMEMfs6JkoTvcezq/6RntCOcD6XYNvovSK/ubBKg9buZSshDveJlrJHV8NcA
OTSLF3EBrhaa5Vq9WYdkNz4zIrL51RXNFFa7X3q5Y6MHeviVhI828uhfXgMdE3RH
0PFu6499DrfuWSxJ/fMkoZGjp9HKk5n3YouZQ0xW0Ir7I3wk6U1S0NSpxLI+ZVU2
mMI7nx44Qtsi5GwCiMgwriCCplVi9zbAwMvbmF+qBy9V3w0ZsuOgpQj0OKkTzk+y
xei3vCSPPLv3oNSz9RR42rc9r5e8qSZONy9fbcFoQjhAsLgNlRBmaIS86Nk1SjFG
FP7/PvSxgfeupJYutPjiY75+zZNS0I9MgMK2Lb9S0bdDBpRqwHIMCF2qbIVIE2T4
UTnXqTVX/wflBSMkINWo4NrlEy3z92eVy44/cTOEY42Gsy2ehw/G4aXS4Ps5jN+Y
GhuBbBIE60ZMCUX9TpkQTaZsdSbTxi7/R/CLRSGF8LQY4sdltezMkoi+WMCdu9Bv
GOYyz4F8XTcuAXerD9ybMFdAKrB8xfohhYivP02lFN19x6bMgXtXre+InTqdivjF
mM5DOOre1+opb1BX+fHozdkHhof5fhGaCJPb9bWrUSViaDfwHirfGUIKGrlfcpXj
th9++AmFnl4UKoJPmntL4IsJeYffVogAfcaIX9BoX7bmBrVSlvS7Rf/63vRagV3u
hr+7xaLULPqsq/QvXOrsNCQ57UCl9XYxVE4rfG+ZDIhCcDs/B2t0aFvZ8TIh5qfk
ZVNqkubolFXQnSTX8vm1/fI38KaPselpSvK0AzuaFp+0uVYtwMHivXWaQScQaAUp
CZTx3fY1hkpqPu9RIzri21Qfegwy1TXVNsVuTKjCSYzUSkpgLh2KI5RUVcvaJHh+
YEQVIw3h5TfBits/HqEMNUe0chttgIXm1jFjOFmJf/UpssTIN9GUj8XubioTwwOp
Jto7Kg2eKwZPbWhttnh9f1wKZXt3vq8ZfzaJy2krk5fK8O3X2095Q+A342TTy71p
QJB4u6dRlv2XOLOhG1emNsQB6jYQgctJJ2/wUeYhH21XFqydlHqMXS0PSTU5ATEs
xIv+ZL5Zcj5NoTMGzmfuZk1tOqCs+krpAmirx7zWvhr/ouP53G/N5n20Vvz0GeO4
tgFS0H39+w29tajPH3chOk0YKz0R5hHFQagDKvZuus7YOhL6Tcq1XeZLNXHhjl5Z
WrkcRaKuJUNS3vSdnuGe8/MYvNDuFAR9mjn2V0gDjGaNYasvIprkTKJM2HooEJtX
AvFJKgu+bk3XDPFjr+K11jqNzoixB/iV8An4IqESBG+PYqjQUQwP5oewcJhADz/y
M+gbA4lJ96LwZQ698wp98XMP8+2sr2my74zdyR+LM+FV6fizZBg899caEj6hiSic
fRMIRWTldx25rYPqIgskIo8aeQPj0uTggx7F+us6wSySVQawXGUUP2Pp0rYCx+lV
cEHzA+gatie0I7lxhbKd8ts1B/YdT6EjgUIwv25OcV1wSmnOtrvU7FSpuTkSOOMD
zvLu82IPFO2XwTih1GoT2FZpsVceOY0cPPRw4oCTT5OURaBuq9KQdmpwm62ewF1x
3cLpFanhdnc7BxJ7ARHj6CkHTaOenZ2xlsvho7GmhK+JnPn5dNQDfieb37D8BQun
7D+HtXLTu2qA9XaJ7Tiy+noEUhgYIR52KyQX3LzGAN63nSUWdIWpaNmCMoGNorw/
AOK4VtBzKDnozbCbh7HyLY66NaY4vUIOYjIAS+nYJ6NNRbcngPcdHBaXylMZ6Yl7
MUiIvgnl45inKIm/OSVpdOCIp5fPBSObboTZ4nVuNC+w8K8Oq9D/bAzToLxCKKRZ
qiK5uqamjQHUngMXnDE2izgO6xKCzapAhsGDz3pFcmThB0h2rdt1MERrOVFYyrFk
HH48tMi9jqhJ+bJAnPAHOnUJ2PzjxDY3RmiBDqxAk4mFN8NqsoOsrWLBKcbf5bcx
izD7RCbhpZQj4IApDdQ66dSmj0CcKgNiFT2FnOXyJ7XRUC2DGwr/GtgF9eJUzBhg
Ga888Su1+4npUQBrV8Sv5dKtkCdjQK+QbOz9hulVgZ1LNTjW+uZF5N2QWy9g/ezC

//pragma protect end_data_block
//pragma protect digest_block
saXiuKN5JqznsDjEA9SSpNGSKdM=
//pragma protect end_digest_block
//pragma protect end_protected
