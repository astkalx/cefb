// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
MW5EgWrwkEBmZljOf0SWSo0N0+vsac2Hb+B+uJQsS5UL6+WKaybGkw0Sg1KNklp6
q19AJDWJ4B4XGwpH93NtSAUP84ToN5mvyGYlYGrG+5NbBEfIQNblmT/+XYUA3ahB
iDZ4WJnoVAQKz5gUbCj0lBfNzNHFFTiiCBkClKRJlRjAvovrXxBbDQ==
//pragma protect end_key_block
//pragma protect digest_block
C8i9PqHkFiA70KTYMtM5K4Xtb5A=
//pragma protect end_digest_block
//pragma protect data_block
2Uj8jFjo7plsaluzQ0CtmZHyXynvw0B2Ec7wpCuwU7i2Lzve19rpLvtI7f6MixLk
h7sOM/3sI8+3ML2yWpVX0Crj3U9bawuJx7VzIPUOSXpYd96Zokulp7qlcyZjzDFc
eQjlZFJ3gmxMzTqoiMD+aK/QSbi44bmiTmZpevw7Dq3oM1dfeVfF36Beybb4dxvw
K8+LVZVu5zHj9XfYy3ZvHQjeVsWFiEr+vmGWofAiE7Ka8X2lpmbhwZah2r9ziBgJ
RocW/feyxeL/AM7Mqk1J2fLQbhpqyqADCBMEuN/KPc/6dBj9NM5IBduKspallh42
HyzD1tys4UpJpzd+aZkheNzlVGA+Rx6SsM6Ew8RIHPTgIrqH9qYZ6YRGUPvjISmD
ODVO6tFQIDDc8vQcM+VUeYwNg7hOczU6SjPraedwRCxI/pa82fef41RVxjfM7lPi
uYzpM2PYVtLe1I9PXhO3I5ajJue3bUaCPVkbWv8KnVctNmrkxDmxkr7Zks+h4JL2
eieiRPD/P18QGG5VICTEBdM9ucs9rhi9l9uRnvtZAK/qqXdR1wpu8/DVEXxfQIOe
/vXseLdD9Fq3bCsSzdxwKSM+od16DEjLECcOG3dq+PosTWEwkYBntDh5muzWrMH+
qfuQxYliv3QMNbi1wTRb1pPTP0C4pIDMyYFgkwJCVGIvTr6am188Zr0GVL5HQG0/
OOXe+h0v8o31yBX3nEfLNRwU3KpYIFcb+SQm7ekq5y4q+okqN4gu3cqjyvALoY+5
BOZ4yRqrPgpI+TYqbd3BXt4PyblTb6U5of0FSmGEj17gELrSJy8LkJgJp8jx/N7g
WM6TWhhPZTr44cWqucFRaDiBpi8nOXdn80aj/KQHkQGrjtmz/Pb/vTk9yuQ4ufWw
Dsbh2FT2ZQf6TPfdVZbDwKD4coeMh7u+3eT/kF8phNdrb5uz+rEVvTzDsEKbfgx+
hm+fIYKqjLEDYG5lU3Ac/L0wWoKUJjxcvEJ4o8j24iWZbuPmKRnKuqziulF8oKmC
GhTePsQRafmBBcZE6G4S7Vk87WfnxCIlP/h1Rr+SLeV/NSJBEIzih0MePZ5aLDam
51nOrY/5OpZd9yunzQ8aO29m3pI7Bnm9eqfJcjbwBoS1/5XxMHW/FpfW2+2U0fWE
eUphG9CqiPbom4THmNyeJ8JzDvOkMMHdeE+rvr4EKuKwc5b5KjiidNi6bSJ3kWGw
6uTl26MpRzXe6HRcBeBuiMFlHosIzQQ/Bt6otqlQ+zsYu6Yc+NYdFIvZ05BylVoo
s/qNVNrgdbK1LmKlGklJtEpWUpSFCfwDT2DKP+RRDP0WAq9PI+KDGl0DkNhM33cR
E10JCjilANfa7+5+nYUDtwRav76IEVQ0ddeXLCd+hCeOV/1VI3U0DYD1mdlWfyxF
uyamAndCio7srRxstuD/fem81oWunVhL8eN0KZ0mpOh4btXw/N3ZkS3XkbA3qcps
ZdXa6/mSHS9j3Ve2fDkgVN4GUiQ3Mj2hibZePhDB6FbuWnqwwifk9D21+2JRpbMM
n8bVv0Dyshhoi5NI0xV+1knv9pHjBYf6N91Wmd4ks0mCwZ0ArBEOWfVQV9X3+gW2
jVvWjAru/MhmCXf8IxsDu205o1chOtcX7qj2f4ErB9Ii2IvpXj7A4dVl+gt6zG4/
GBVG4s75eazsuuZ0RX/BZStA8Y2grS+3CBTq9wH5mNbzTgzKokIEwN75LK59I7yn
TsydxNbkMNcX20DvMsEFPv4wKNtoZ9EL3UsVwAiy/nIjhKVGkVxoPnrA5fbuWTcS
YZDOeapGYckUGccNqO+gNwoc8WQcMtFg6viIrMPAhrqsIfcHyeiMDeHC6gL9Zfnm
Y0oIrdGaGfKkd4vTTmjdLAEAM0lJu7EIKbgjelTfVLygPC7/l13vsxKZG6lL3yZB
/R7rvLd9Wu/aXoEeY6o4TtPc9iu+OwxlnxledLHrEULLC+3RJx+QOOt/yzaV47Du
2Y0clXT8kmJF5j7rgtRv8JWC0J3lUYKQBksKSkDKn8Dt8yBDjOEr4uJmGkZbRxKN
ljqFaCHZSLobGnzrSKRXcScMVql6Tcmj+hs2x6e4dAuje6GTrv6Nl4ykqniccto+
EHBy+xaHTEm8NZpwWGYLfNZd3lXdOoWwWl9o8qVl4IWsoN6MqdxWFg2zcoHwFZQB
93FZb8HEE+Jhxgr+R0nskPyPIC1LF2th4LaGHqXJ5Pf8nSATLYxXrW3JzQDYGe31
/MlPZKbx+wc/Zzj1NoVNCo3J8+Tz277wgZvKku0SWSSKDFiGvBJl6bOCWwR97ejM
BmbLBYFrG6WUTnpax94ZLVNFAguNZlb8JmuYnKUGiOWlbSpQv573sf/trPaKuu35
QALVKgKDwpyJ60qGG2+SE3yea8CTwo5yWUK6llPZA8coS9zlkTOwnEqUN4M+97FX
DEzIKJ6hYggV8s83iM2A56W8rAHtx/qm39LJ/RrH2vWQVzIihO0uwBAhS4rSFbJX
G3cU0/lXgG8/yiSU3Ysl3cPH2XnQSDn+CLhLejx/d8ngudXoUO1kRi7y9mOFEcVc
1rBMFnouqkPoZEERLTqkvdMeOkVq8bYwT+9QNMsxBvCEaPiTF/V+pP9iYOQ5stUL
z69zNvx/FqKcn7BsAcMp86j+QIfBLgwxUh8PUZvmmXvHX9zOKqoBIGWb1m2WBfMK
YGbw9zEziwuescuB7ZNV9+BZMT5ZIZd11dBGGAxH3H4SE6CcOWS6fhHy0FBl57NR
SW2v+2PARL7N/0LCB/GMuF5hm37+k+gaJnuNfKLAdUv1PdQFC4web4FpAvSF4eqR
u0zgty57bjJ/OUbTND/uGVj5FtkQAK1SxaGsYjORV8ZJdvxqro1cH2Az+xKElK62
obL5B8YJXyhOa+g+8u/9fRKGKzCJiZTCVXCukbwEJAfxHwliRR8V/GnUDg+He7Zb
3RfEzWZH9NO9Ayni+KJYkpdOThxYyJusDSCTs7uAkcC+hnD4KpOfwgRtAEzR7owH
sFWcPhfGQDzvCG2bgtKr8ByTHfNEWPJaqRIria125YY4U7VWy90kQ7UOrT9QGXdZ
OBkFP0jJ8ME01CRilfW9MDrHJVnXLQOuTqJH9ucJ3q6C88Xpez4jcX/76VSpQEXu
8AP8Cc6iYWiafZhCVm9bZfXzD3Xpy35WLqcofMsaFb16HmnfNeG0Zqy3gdDdG5Ys
ehcjDXl6RD31hLLGIW7/Q2d4ls/jmBieksATBNGW6DKXZV9wG0inR11tXCysWD3p
QNKjoyOAH9Ovwmd0u07at3Dv/n3fc3pIcNQVfnIKcpqOGLbcVgKO3min7d5dy/5L
DEslYKlMaRUtKgn4ESqfgMwq9hFZj4tWiuIpDSokDkbQ/kCqz9WJbgA5Lxgs4flN
QW9PwjqZCbJR2bSXebKPqhbrGIDvBiQd6Zr2QIFK8yXb8+PxrTWisYLftVPCnKkm
r8OO+S7/2ldn3cGXbgnMPckGMLdVOIZdr5ayYDyA8kppq64XJxbZMXuUfiFb/Pys
TZbDI5KHakxYISZoB0oqpjmmmqt8czTFsoG0iO+gJ1oXIT6MqZntvpWO89pKzXhH
UBfGVZtfm3OhERD/ZLIUhe6/gJNXyqiTg0OG4XNgvIjKe/cBx21jm0GahS3NOJYh
QSTz/t2911MNB9q2uMCt4G4m+XcEgvNiKhOZllECueBlBmMH41VqXgZc4YbJMSV3
k9jHIuhWeYQTIM/emvM4rL/bvAgAhLAiXaX47RUV6SmsUaiBdFchySMylrwVmwJi
lbphM9+h+KJ1hZ4hGsG9GLmuKGkzxE5WKrepeARUHhNiyqgiR5Kmsh4OyiQVD5ov
0auTIlbZLo+PWVkBEqhwJ6CbRE9w1DVexfvpfCTpG7cLb3xmDXBlRg7vmaFvKjyZ
I7Z/sLaUU5KOCCaH3WGHG+Mn1+hbVatGu/IT6w4ebmGrEW7QcTEIv4DCd1uEQWYx
LK/1HAwHvOPbDqCSvH/HoVd4xIB6EQGyxEgmujuXaHDSSgotl3+dLavMbZRAWXE3
dS+Fm02utncB+eMqYJp/Nv+ZJwtAbDqNfASxqYE9RP4pwnFXC+hKGH4DM7R+OWoe
V74HrfRtIWs4hX7vArrMVWI8nUFCewWOXG4EO8dSj5OGJ5/0KabIFegxxmxWd9Hr
DKOmodzjKQhlYyVxPvo+bV3tF4JWSPFFrML8tGQ4yNMVONt+7+mv8Hd7ZWJf0NNb
a4Gs0yCArewOou361xDDFO0nq18g4KAuppVFTGUSZzjpM1G1F8rICg7NdU+MXG23
2Y0SWLYJEVTEAv7HjSis8rkWURf8UAOPJNZxqhaYWp42Pz0u7damlLxvXmIn+P9O
VHW1dDXtQYGJNutitsl0Otme9Dkr91x8vKXS0c9zxLE+zQyTGNmmwGijaa0sGiDr
gha0L/bpBuT3LdD5lztUOnpiMiPXmtFtBWLnLvqtVg2nm8GGahj5StPFTfQHywGe
EQAqdnsLGcPrFkHMY8+W5jmXfpsRF1HKdl+tHQhK8Z+R5dz/0ifZcGcOTA9aDj+v
eMlgot5SywmHydOV1I+fMAO2gkkf5u63E4wL+JEOsuYE2gjgcbQUoGwDVr/7dOQ+
OjIM0BFUOHWjwnLdkrrGrjWSN+iGnsPjzPZs8S3OcwsW78fGQdko8cIlwqbXQ7p0
J7Cu0/qT40vlGrJPuXTz9f2AremqxMyh2L07fA/v368zbNW2rjGX+D0TDhS2lWtp
4G/ORq+xicrscUjSYz9nx7xB8YeiRLSpJpd0PpWhtPyh4AnBBsmCQeCW2D74rmky
faphOtAREQRYH8NKXWZ8PisDlTGXVpSqKZGVkLR/4vNZF/4nOJjkUdzs69OI6IKK
NO+9uXW7iM9YZINw4EYSkDf9x9yNcQnPMT/xbopkjxI07qO0Gu9r9xPiwmhXBWZh
FOSnplYLNTLwto/IdVfxZXPKQoz6qBNdV6oW7x6xyqoPwPj+qpA3V9rv1Uf+JQ3z
R3RjUnDDpXRjtJazBqgtwOZeC0Rb4LeYSRL0M7FSs9ghnVj5BFmjJurqdhoSN+gd
r/LOHLolxTSBnaJspBp8FLCt+ciyPZ0oAMoDt1wqsnGsjpi1u+rsbtofbEWUHNFM
cj7JA2quUgW1C+8nYLmMZmHIADASmSqKb00VRzX2ekdAB0f+IBIoMsQVttqnNvvE
KezgfbdieoLEOGuJc3ldWaB/ZU0ZqprTNHdETiceDXSadO0W7vI/A0MEPcxnOF0V
Va1x2R/Pp7KMdIRk+ZLOmtuADpy1lt0xjoeUMHqovb+ZXxF7ShEVnYqrMjhd8asH
B3FIFZJKSfHtTETAepmthp60k+1VJCX2Ve34s1gy+T5oCzRCEehF1/A3Zt28xVuQ
ATG8uo3J+ru5wbelbfqcfrFm22F0mOefTGQZKjbQ+ghEcP1rVtc+CGmwy/LknzsF
65cOeDVFuBFxo5/BFRzZgMXmyvwKAOSgfiygHBIjSSgWv/m/+LuMgH907s/fl8zl
IljFOaGnEWKk3ZC40FhOM6QgW/te8UeK8gJwpNHa8WoCmEYSD9QRT96qdP0EOqI5
cn6VcLgo7fXAbuo9VeCXIktl/du5qWOO3LR5CXsIcnOQpD9WxdKd/12GS3+haDmp
2RQLUfZjZSoU4lk50AwNJItS+R5tuMBko9J0KslXYfGiumFZHSA/h2XfUjbsqDJ7
pDx5yRW3c3QsjFr+J11RR8zi43VytlEzQokQdfr/Q+AyzifExYIOT8ntQQRNNfz7
8dZ9iH4bKzHT1eI1suCEKXLjom4Wg174aRIPScZdGyEm3CmfQLoOi02zAcNbg8qD
/D+2U+FJAXKMHEi5Pzs0LfBQIO8LPAv6R4prhzJ7V6o2ycuXCBkaMD6AJ/vvDwKh
8CPcMEbJj/6YAZ9xhfHyhJKch4KP7MScBeS37eZLkA5eaNjfFASb2VpYK3OrpYWG
b4hyoM4V39/BxnIcanQv7+WKw9Mt7GwREPkYXvslsmjfNL9l7qbVIzidHLaKbRkT
Ni3JeXGYmupKOy0eO3yI2pMrANIZ3aSDqdzcg4WQgCKFhDAIZwP2tGrWJUbpazvl
WmeCfuG4A7YMdalQoIPQYrKK/8Za/LeKT0peI4nSJwr2iRhprnBY5LsfGju2dVmh
16vlCLNoTi9ysyLo0jRTs3UYdXDo1ibI5HbhlC4djAuRPgRY/hQ19uYtrM/TuX/m
lgqE6RCQDhP9LeX2cWzkBhg2GtZpu9VIE1S3uVq3GPWetTiXynD5VehSWthSH6ah
koSpzfO7bFQ+2jExK4SQBKkxrPa867/zP9l7b2nu3WbwCaHspvmRk7YbRZ5hj9m8
SDwoKkVtDn5BjgykkJh5i0QF7+jx+ff79PKvjt90jQ053oqeFBz2i/PlN3UO4tm7
y/efKcNoGkU6JtvTuFt9xLyKd/dCp9WbA0Q2DRz2hhzP4/DJ07zVsvWzlZ+a+V50
PGRvnxY29USNpzFQYik+dIzRKNxz+tQ2wuThNpMU+RPcrbehu1mwUNcMBzfHZNpm
KlUsLr95uOwMqI1dXKx9S6auOvwEhMQbOI7df7FUPqrLByMEtiT2KwlySAJxh0wN
l00jY3N6AfxLXrxcM3K/NcMgZLHfawLUroFPcRo0Mcu6NSOTh9u9vTT0cKFgZKOm
W/14J5jm95zKbPDWJYynygNXlAA3gadbF8/NXLCXsRpXp/h5uUKhGheurrvLmhBs
WORM1qPYPmlRPvlQwtCYZ/fyoyeJuxbKQMmF+H6NzQrQscBc1f6iVTVj6VyUAPKa
gzbskPLxMruRyy1jzMsLD+2+vsx2A7lSRdBmwg7O1l+zuMtw2vEq1R8Ly8X6Vjin
87xhWYHjznCxb6FLtTKCMESDXo3Sr0dNHqb9QfxfVw0vnQ8cV2NJkvcasUD61oBS
Rwlb/Q5iqfmEfjZdaPc+yWMww56CPNCh7UFfuQ5fcDuTfH1c0XkYiMwlgIjBOZEH
cZRMpmLaRobn5HLbpyNoOPEvOD7Xg1n4rfpOBLmrjZ7gvJo/VdlaCUh9qI3oGYTy
SBP4YOeKcK2ftwTe+XbxsApxmfc63RrDhnkCvJyakcPHh8r+a9z8pvKxXHPxP7rd
tH+ajrTFwYq8AxOMoBai6M90dYOnKBkdJR+n928Q6xyoIBz5asvTf9LlQPrN+a9I
/1eryJCYcSy7hgZc2UuujlPDe7P7RuS7sFpfWsb2j4WuTvmmvvPgLJWXgMbc/oLY
e/i5KonkwDrL+8faUWB6kSdY5xicyoJyVdJRqdHWulWqVGqCMbK0QguoBrGGqRpu
UQ4kqtUr5pGg2T9UPpEBCNnUsRwlz3bU90jVMrgbjUAYMyPqwf0VPix6Cf69yyEe
hrWbVETD/R8wtUEXKI0txUJYWEgPV+Bzsar0dgQG0MtQKhC6vtD1jjkGNsCpquZQ
9bgQipyOEZkFFOgQ3ZHb5fjjbQUpE+5xhIz2j65ZPuAIREMqpVwpzdvtfGS1JV/0
3kCWQQnl1kjrsRTXphl+HT8oIKhQKFoDlbPZkhbUhK6cMrr/5+CXllhTdb/v1OE0
5mgUfx5TlhB0KAVVTtKPCZ849RECvVyOZSCim7G0FPGM6PbqSpFS/riWy8QtjRMW
q2kfR4lm1Ay7Zehv0S7KJ78DjTzwPntX3FIhizrueAyYjAd8wMIul/ymcNzdrG6w
RGJWU2Xz+MS9KRUiP+UtYDLQ2NkbSsZZCxRheeiTRRpOZDR11qV6ByMYYaIFvrZV
Q2SSQbogJPGaUZ5/dXB8nhzBxrp4RNRtwpfXajsm+4M=
//pragma protect end_data_block
//pragma protect digest_block
v8Pz2WvGsqj6zdYdtrBAWyQn7XU=
//pragma protect end_digest_block
//pragma protect end_protected
