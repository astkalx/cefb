// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 03:42:18 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
liwEV3CLWh6CC+UQQ9wH30YNBq2jWySuB1aMSwbxW1XhroJrwaoiEbrRIOgBz3ou
S88VQBdKqYtzHh+9u7aBz6bahW812K50p4SmTtmcAZOib7OoK5ZgCCC+lR1nwTrb
GK22F1hF1kknz8dv6jeyXvWO95/aT2GERykj1eIWPpY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5696)
ScFLhTZwijTYJodFyGssP/DRzVGfi3VnuBrWYleK+8z0FAy7+lbFrfNkoUEdGT3h
jc/WE0QeckrnY8NKGMD0IV9YEs7wuOIOWYLndl1ge9ivQ+GMsxGz31ZW5CdzJ1sL
iBm95UjDHiRIoFEtdkrq6rrtNx9hkMQeIXMAdZwqOtTYjp4AXzxj/xV4ba48cqfG
m+cx9Zpm4flLAIS6V3PXoUtBwQtA539CnEZxcTrU4HJ4s5kB9nslRdqLewipkBiM
IhDXozscApe98opVoMZL6+Ngx9bKVsbc5gdxbKoW4Mbs9m7fIc2lTu/1Vfc6nn4q
GjGq8wAgA+zHOUoeS7r/qDr4xUdweQ0l+yycw/prmkYrev491fGgrxgFINF0dX/V
ZpZPFeJQJJhAjOWniMhL0ultgt4AM2fMXzyPAHc0N+s+NkCFAqDHgH/mfrv5vecg
NpYv1sgxpnynR1SzMrE/xBC2B3y2reEaZCxEPyiQFSxAeJzr2fBUgkWeUIMLEZw3
Gg0TQQ6VFKTWMk9hqA+w8hTjzocvJgH3rZYWQBQGUPkgESC8aJCSVgF/ge+3wpSD
kc5B3xB+S/9Rz2efUBwVLpPwt7IAdUGyzeoeV7x+UoGI/j5beQgRmwCrmL/bKGJ1
1JtbF8SKHqqSXREkes/WhiEAjJh7VCfZvBK2T0P6EUrW7vxaQwCZIckIuQNy5w8X
CV442oWmu8/QGYIX/IVHm9sulNaPddSEYdpU0PnoT3fwP89hIg6ygWogXxf+RLcQ
SWDkL7HTshgbzG69iYynYX1vKUnEgeKpwqwXL6Te41FJuw9LXHnfGmH17yBBtAgV
UNOjby+PBoTr3nyZ5+BjobLyux+nCrEVxL7PqlUJhIafSwIgTzYWNiIH80vaJXju
BldiwuzjxusqgIX/Pww62e0ITSTcUE4WjUbtBeDssM5d5GX3YnomRiW/d+ypvAAc
b9uVSlt4Q2nVAyeZESBhD6udkHDC5DlPfGXK6tEKCqLyLUjAGMpweZpycBGN9MkI
VTgrnvXFY6dxwmGksdpZ1Kb521G3BAovmASEcQkEyScJnbOt+Va42jBEWNMjqKsZ
KtM1GemKRph5henSi9siMYBmLnh/M8mndWZKsdLr3/rU4C0YIN/w8W6pnZdCeoIY
QVynn2ISNzwVz4eG8Ak8azCg1PYYwC1SS5FaOILo1ytW6pKf7RdOCE5ToM9Tbs7a
2XllniAX6OWD87SNZH/y6fheo9LFVe3bDfnWZojJaevXa35woy8s6y1k9LBL0YKJ
CWy78KSiwc0XV0oAn6I6VVkDqnYVHeKA1vWTDzCqaYOj6kd2l4k7joD3hKw+4G6W
XL/cKmRiLpq1s/1QYzLAJfdfYAHD0o/GyOrxsCgTPSFeYO+g0qqQOXZTT1V/LGZu
pLuFly+19UopbTsFPeTB/PEXLOihEwOPvM28dALNRqRm9FecttYXGJrUvlgkRdTm
9QX83zNE4e4lB/H5e6BovZRXQfm8Ge2Bt3LIuOn2xP0Tlwq7soJG37akHZQMwf4b
B1ikypf9LHBb0gQuG9U0SsqC4YjEvtsbRNwWzBQztthev0R2XT0j/x+vif22NA+A
9enjKLklKILy3LGmh7/2ZPbtIhhuA4z9Wgr8/p++LvXUN7/CfdZGzYEfv3ZTS04+
VaPeSDRu4ZEeup/w5+n/S0qH3GHdticxA4DABqLD3zKtQt0NgE2fkRZ4zzWVeQdK
V9t8cOYzNf7w4WRBhkippJrD2pDHDIC9DnvLxTGFXIK2w6xh/p/dV2yQzAJZl+kp
lv4xeMYuFmKh0w6rOCD01CvuZxGWAFEdZKpI3QV9cb0z+vyVYn/e2E7Xj9uqxR1g
GXdvqiU6OvYxutgLY/iW46bGNva0tO6K44dfEwWMDlfrQX2nxNluYLHvXJxsWGq9
3jpVa/VocRssyoR3T1rtjoETYO1OT0eTC4GmBzk3z1b0ES2JO8HVCrhAhE5dudrP
A0N9ZywVxrUw7oVPhTJmE1JrXd/bKhtLEJIM3sa6/+LhJsVOsJ+nzmLK/afQGQiH
iQemAUdHkpA7klCnDJ4qssbgQA2W9I68TmZrXajUcIpfygYPgvNt7SvRYI9f1PQl
mjIIITj6M+h/xSg3DCg1fsss0XmgZvpmVVtKtTwM/ypWZWjWO6Pz4q+2QwHB310B
1QRKYq7Sh9wmEybRsT1wu8jD4+/2D1DCdkS4UPQR9pJ2uPfnjeLdJJKSlJXRJwVh
dI7i0QtrkI4LuSuWeLMVs7gWtbeNcVdmVCgIHBECp50GrLmWsayn6/oSvCSTWU1q
LAm7xnabiU+InhIPp9Y+HDPAI6yATwY2hNd8jorAi+TXgDkizqqn0qQryfR+hkMx
OoTowTMAuSM/i+YCqymUwA9PBpJ/8rEvxvo7HwltJ1fe8R8Vpstp6XZ1HUpkMh1P
H0O8q5Vc29ULkkGDReaHrHj0vj45vJDdAKhticv8UvAYp7+BLb/THdM6looaHY4M
EJaNmZQ8tsFFsgizqZx1Rvxwv+I3DgHwPMOx/E43uyjZIPXDA9GBHQACwdb6QwJA
h0Hhu8CEcPeuYYuxW+sviZjskYjOVfYcE8UqIHp25ZS0pn8w0bCvsolxdQw/OpCX
IMgZQAa7sI6INUyD0v1IBfMQv9CO/KK7nmWS4g0UP2LEya1ILdvSRKsjY6KDGwkh
CKW+LjLpcKomKdJKSHxEu0rH7/8HSNMjDIhHczIotFN0xmrF7dWoRB5KV1hti2BA
kBITWE10MCB4q2vt6NfRk1kfsebp05F6qkVQlThV0uYZ+BsC4bt6Vj0Fk2l87/n5
rfIzVVGbqfm5VKoKfiXMPmwgx55IFJoP4+l/X7Lx2nMEi5ZJMm/DY7A5bRto/lgP
NoNdjG6zbXYHISSbRMDuODRvz2d3CmuD9kO8TFPqA9+eyCoFI0DonyF+jFPbWkP7
sGlDKwLdHbSmd1WRcY5EdFyX1nS/dZgU7XoIvQXQhwqJA4HyAZQ/2CnyBIdvqG5j
dSnOQgI4JkQyeTeu429epAUKKX5ej3/YvzqH1G/BN2fZlcRp2ZsWEUcNNj2waKwN
JRwV3LGenZFb7YfKieifth4WhHXNgc+ojHOodWD3k9KKbP7XjbIN9JJkbu5tg67P
MYEowJHmsQwPxlPyk91nBLmK5EAB2691RK8vAkcj5g2bzbKBOXyETKBcLzEJUxnx
qXBGKPa3Y3W9M+1+wT1jdCeXF7CVvmsNm1sl3rXAohr3pLvKtEUJCQ1El2eTNq8d
5ddSDO2vBnXxOJ7IAC7E9Z97c7jOOBd/RG2R6/yXRHgkSaLe4eDylNXL/by9KO/U
hH+MWQD2ZBW+GiIO/Hlbt+o2alff/ViSsUDcMXrUbEOoewGFsOJlIz9A4gqFxrp5
s8b6sguFAGaM9nyc0PNf3R+PbFNhkRXZXd4iIv4zutBNansEyIcniYeZgK3XRnRO
YkXb4ElEKun36mqqCdt1JUnVizdM6BMHF6IyBgIM0vg9yr4lRJAMl/dBWpPJoS6h
hTky8OSF2H8vrplvb7hFIvglh6V12CHTx+c4gqFdrg1q1R16OlpDahJjkBN32FzN
lKojTg61/7cPlTTWbfqQiWxdZN/E2gFCo0VibZar1xz24wZbYIGsV8kY1ROToam6
U4GBHzCQz5DlBujU3UcP1mIn9ESigKfUx3gJlqdbuzvQVS5Yka+XrfnDYFZYWD7f
g2Gt4lFv/HIQ3LJ9WTNPntdYus4TPME/O16+LiyRy1SqT0FbaDP7t3CvmF7wgPmN
HWOWHiHz1KOjqFuvJDuhVsmiP4MAr6+GT3up0R+RTSKM651cYwGLMh2ujz9+RQDm
a5ufXAqbVtWuk7TjrL4Jmanj3Ft0Z5JxgbO2REhO1o/pcKIHbWWRg0QNd5JgA+b7
4pLVbz3uLb7U7jRP//esJ9ByMY50NGsGiiyyPGSmKrKRXOKtkWDX2ahJI3TW+h6z
H51M3zG8KZvFbR8GTX6FpHZvWoRCxFKsupahwNsIA3hmZwHSLTeF7qUuH+E7KZFx
4cvt92WIOJh0ueAZ6csE3YROt4VqfGn+802YCZOSEkVNYYf454uZktCee0VFj5fC
wVZX8T3rS8csArzDgniaROvoyfpTRL2tkzY/uJQsV+EnFkw/+gXTNQ/yZpiPJDED
BPQGdBgrZef04gOtjg7TftNdjmPQg8xg+qAIb5gMGlQxj670DvD1+dL5XePYgDOs
ATjzYd0NvcQhm4VQ/eDjQ4vCi5JliRjwchtQhcJk26Q0l/r5ibMrd3692DmKX2be
eKk8ln4UbOamuZprI9WIyZpja5oRGomEb8nsrk2jQRlE8Jf8vvNqMCejOBAgl5X5
WtKv8abEWBd47UeWGENSNRzzUhiIPBlopNpZkoiSONL4DkDIVEmm24J120DhrmUq
sQIAylcjdOmAcZme74x4SVU20oZFX5QGOMIbk9XqhZzWx2CxtkfJm2+sP/L3RrbD
eRitp/bfhI2hNyjIRhAgxX2JcjPiXQ/VHXLGthNYdYdQgX9PDp7wtZL4PzSkXzdq
KLVfRAWBzo+f7boiR63+Te3hNyx96o2QLAYyago6Lqw5sABWoyGXDheXH12sfiC5
eiZaJLYcNg+sWIxo31oEvefcEVgC4LXoNfx3CqB7EyocxwoMiSZL+tjmxhy3dbHd
n4YHO4ZBgrh7PSs2PsJqHBHEi76eimfyXWt/CzHa3qi545V5h2hEISXfMS23oHMI
Fu1fkgOHB5OfJHzqlYAK9G7iWoyFplMxFEu9zlQThN/OnDrBjOHGTpSoDaQUdOUL
F38Za/2gWCWAl0CF5SuEztTEgVHvlsrLMtrTgq+4QHf95lm1KMVQc31U72qrsDw8
jEfUMBs7IL718tzX4acvkZFm5wHJ5PPMc4Rk3zZS93KRJIEMYthIUXnyv/s8mN3g
6jNcLK8Hxgh6milKiVZ3SNmxYtT+W/QBCwPYWhA4cJWxFSZfI1OyEdUh1khqaVlU
SoBVMOFSNyqWosmxqRjBXp+m1bHoa94ovcXi0Q7mqOE+2ydgXPXhrVmnh7Q2girq
d7jMq7DJODsDLOdw35uuRlm2xlWTjO4Qg3H8/hHzBEADCpziAw7AKXOsmBzUPI/a
tQ/3cx0s6GnJO8AZZpgI7dPr5yeswr2TlQiB+J4rV7kQeBL1AJaXEHASaO/qqxwG
JeAQ+gkf78xlHtP0s26pQv2Kngp6c8a51UbC6STjBXj5Eil/xkq9iUPpVl+eVsMT
SLcbP8h7p/yO7gFyfPJVFNYooLydo7DGFJ8l49dGrpdJP1CqpMlFUJrXhExO1n0o
VRPR78lTbydCcKNm7CPMy5i9sweVpCYZJxofwuMFJfdjFdfGifyck6q9rynRX+lU
YB5THHBjONvZnJAvB1/sMjLPcYEmtHBeA52DoFQBCyx1ngs3ahml9uJXwSTZOg7N
Hl/1Td6locQZCB+tKnvhzf1vtzZqyI4BiZpKSk1UD4pWt2R34MPv89Ey0pA4k0cq
19oDw207nJFdLCbyihAN9LcF1TAlJHNNHWY4ikuFXgQ5T81tpt0/CdITYeuNt5hO
BIpd7svqFM2BBupinJaneX+cLS2j7v+963fIaap00KSw6RZZ8BkWLWbiJoQChILg
bjMzwiiD5jz9hW45gLwGgSp6kZiFOd9Cndvi8T/fboqROAVSTLbGCn34W3qS7tAP
mjhzQgxPdYm7yRfm3dBGC2V6MVSEutIb+hVBNgpPrEem2x3USoOsydn1rqUq4hjU
f4G/2WXmTlm8sw73nfLAcQ9Xw1vjeITeEJ3WZ9DF7nXphekADel7WRCb7WwyQUDy
CabZTJu260rRY4mK3qF+b1Z8kQXWXNPxT6aUF78up3a6sYqV1tiTaWM7vP9t2DCv
kT7jn/tcocy7r1LMkj6QNr1QvxYXGqgGh6iABliuZPmbF32ThorkYhXnCHWkC4L7
oZ5NV+f7Hx2lCjN3blArOMHUeN4B8HqnSeZLMhLVnPRIy1+bINdS7r1/wJpKu+zy
PjsV/1NvS6NSmL7MP8OMtHFlHB6ep2oClKZXPQZCuwV5QtcZ2xBU1tBnF396pfJo
hnL3tebDIF7h73lmU9UlCRyY84IKCaLav9J5RCFWePR8Cvk61d5MF98otzZQe30k
2VfqwH+XXH/wbaGHPBVqyHsqZ7oBl77sx6BxsrIGPQ49AAUJ7gwnrUHUreFo7002
rQedll8oPfqDnQsXd7z1iI19ur9Ailw4kJbnkYsKgtRVpdjKaKnye1o2VrP2cTdU
e5LQ2Ne8wClvJVp6hk9TX4XtHiPY7XyH7CWHxqGugI9Bex59wEvKXKQTwTrg3sfa
db9t8XhTmXCC2ECK4zOjUkTIpFbarz4UnPnplTGc/laMTezIUF6Xk2dht9yciukZ
vqJ9lkHvGyEo2KWyxiHzdqJnbEzhdef4NN1FHS3AEfuF+jRx4GPGeMXTUTEhkGIs
NVedInXZI5qBKjdiDLLHicJM8RUfPDEP12qvHGG0g7mRcT8+ruVoLx+c539+T11P
dcj2r/IDwoa+34EmRGejkyHJykVs97Cb7YbrYD1NYnk84ozHRX3CvHoDiltJ3s0N
cSBWuVsQLhjg886plCfFpZ4yEuzAn8wqeArIEbOUv58q/7RREmY7iYbcKSVFrYTz
7huwzhlEa0KLvmCP2EKlm9NlBbVx0FPibFp1ktgNwO+khyQdE5S3YPblMeRmwebr
naWZCbYr+pH3PS6Mfs0HYxqpdsDINbjeDKcl7b5qjSLoy+ifCHt/afy9guvvD8B3
vaJ08FQtfuHd7KkiobMGUIBVy4L5dMax70oJu5/lV3m+LSczdqcE/GmekGCcpdzE
3rmHCZnbY3gEgTZvXCP34fFE2r38yvaiTRqdMm4zIVtPyQluo8POT15LJwSXFo/G
2BjcHYuJUQQngd1t9yG2rWHQx2p7MBHVrZ/lIgVl9mqVXIfhw+vnUFrvUwicb8Cz
HIut/Tfj3Q5mIi45B+dkE3JdISPL0MbXXDsKjeTeHuUEf6FygdYufHs/I5n0oMuY
8lv9bBzM3VQ4MjmWa1vwEOs0SwtPbKW7/fl7m4raTrOjpsETjvHRLd9mvNI7Pst3
ITos4bunpfDDnvlQ/MJx08kDas2h0xtNRlLnaZ/3L1jmebnuwzrq2l4lDQ527W5Q
LDQPHOZr9XlwgIIHd5Xc6Xq2a2sU68ZIV+U7XJK6p6wfpdFwNSE9LfOW4fDwUo7Q
Dx6Wt7wkkuPU2kULQt3tM6A5jV4VCbVI6kHa1wkcyonkjhYC8ikQV6lkg8WzhlWD
Rhg1Fk71iRpUrSwabVrFzAK4KJkNjKSPHVKkCc/JcugzsdZ6SwQWbVShUv3vyd7E
w6T2hASU9y8hQL0JezfiZp0YY0P5xWuudM+LbiZyzZSVk7Rvrh/NYNXxH5yJZZh7
SpK1w+y3oA+P598DaACG/qyzCnasrWaQ9O2JCEdBVDBU9GVYXdoecNymGE2za9Jh
bmqlNLWP5HNnaIsbiE+wF0LV4opneKwZHaC/cPlpFf0Z5/AEkujs1tQ/QB5id9Ja
1hs2kQkKsBGFcIn25Xjc7vTIzwhXmjB6Yrhrdz960UY=
`pragma protect end_protected
