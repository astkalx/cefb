// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
HNPG/JU$LD(+"G(ID+L7?[NB74;5*]^.!;%PWNRM-EXT A"A.41:=]   
HAS@B((*_4FX*P6)?-/\9T*'0HTG,BTA<Q3\^J1OE>G.\>R;DG_<Q+@  
H: ]RZ,=EG,]M<POFSSZM=R@*82Q]=Z6_=[\==\THO1 J^\GMI=C(D0  
HQ02Q#<.%D5L6FYN'FUN/$VCGLNV[>5U-Z[#5KLKK+D_YB%KR\T5<A   
H_D37U,Q]ENQXYQH[\MW)41CQOO8K8X%5ZC?G>=783WB@.,9ZQ.OANP  
`pragma protect encoding=(enctype="uuencode",bytes=3728        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@(2"O'!'U/%$HC@N48QJE]Y-\=VX0JN4#R)[HJ(; C4L 
@F^;19^0-]O2MO;(6;)_74KJ=2+Y!GLX^B542H&:3NN@ 
@O$.O24S!F+3YHH"G@^F7$MO+0*[L9\& 8F\]QCT[0/( 
@"MC4O#Q.MM?*"-'0<K?36UP53'-&GSC8>[\X:)F/*ZL 
@F[)OH%-2,M?(##<SQ>R)V1*6_M<P':(0\I)3KD8"S.8 
@&F,G=3S@_:5!<4[?V8F7]^A&D)/EWQ*&^PY5A!%GO"@ 
@,#AZ+8A< UD!\^ZZ&"ETO=XNZ%GR$^"+<(/WX3\;!*D 
@H%\EQSNB6%2LVO([0O3O#L5V=*J,U'OEQB= 1;:=%,< 
@Q[AN4UC4B%9:1D0(L?AZ_.Y'\4GGY6]6UC@M?3HX1WX 
@:*31MM,PK #7? )?PZS++KY(JPQ-!B&U"[8:^^8BT=0 
@-^@230@3TC%PE#4:#?RN:SSSIEG!;&*Y=5;F4?7$JYX 
@I>TU'K?RE(AY;YU$$^A^PWKV%^BD'X LESA=@.=)PBX 
@)*&"KW:=J(H_CMS.]):W*7*+B3/>9Z SLL11RL<V*[$ 
@L\S=']__1#D6<)&^*X1VE$R,S;9X"X6/$W^HB%QNUS0 
@3^[K>L3?>PT9C0D<D *@U:M1P'XYT[!Q3[%X@;^SK^, 
@M+5Y#ZK]-K_ B4W(M^*%Z/N@'KC<61S>=Y*.R >FT#( 
@2O6C1&S7;,#2L*W]$\G[5?V875P4.+(;7TB@R #>%>0 
@],-E<@96DU%4_,=BK?ZD_X1U/Z?W67-&(-KT+ Z.?'T 
@]II].[11EBN=A@[1P'G]G"C/F^U+^?)@%.'I^]9MJB\ 
@K$TJ5L .[.I#?:/E5,3N^<*HO:WYC4.-?B54;6Y "-, 
@4LG<?!\^:6[E<1C:T)2*_/N(<+S:R==[E]<,VW^>MG  
@ @O8L&QKJB1%!OHP9$'*=WZ@=,FD52I,N@R2W5V!K=L 
@Z>"&3)!0Q%X%"D_#W'T4%,:_XW4!-,=2D%F!/US-OU0 
@(6[8G9?&F>XT M_QP1A"&#I[?R#K\D@U'DL0].P@][0 
@<+-=.L'*+>_>6(4=4_[5"X'X#23V CKCT*T6"4_AP8X 
@NE=D!Y-S](NDE#S<9.*-4"8M7NV\M^\NU2PO8!=3O]H 
@ 873M:>MT@Q<[RBL"M =3,-0KV*E$JC/GRU@8AQ_A6X 
@FZ8_6:-X*^4"16.O=J)5R7&&W<4?RW%7"S#Y^ OQ=:\ 
@1-I9KXWK6_;(3C&'T7@<JVGP8A+A 1.%: J=EB4BX0X 
@@M3>KDVI:%*.4(ZQ19.<!L:%=^HE.$7WMWO\!(XF42\ 
@TY)>2#W"Q%&07]",$$M(B]Q1D"D2)US>$'= M0!#SJ8 
@(FS2!G(^D6RK2GO/%-3$ L@+ AG+O>T$Z%?;'5RC!04 
@%J4W5--U/ J(O\H3*<__]7Z%P:,QT'Q-6O\"*.FN[W, 
@4*CHHBM89Z<XXS:3*]0MMJW4:[ >12QDAJ*>#O:B"=8 
@N@WX-AEYY0_N^WX8Y08*!^1(/C!-U=<7RHDN"WJ(^-$ 
@L\FGSX,],%K<]C8F;W,.E(AQU B>#E"!3-O9J_HY#RP 
@-;N] ?@2YJ/@6#J;E^V34":)<K4',L151"3B^[@D6?< 
@Q(<7Y&P!DY53PYW%BT\1N4\%BP3VP?F&;V0[Y:M8L<0 
@]8>*AD!)TSM2![KD^.<UR?)7V,YSDSAP/Z\;2C >9C4 
@TAZ#?ZE%.,?\'0"?=T_Q5D-(JU\.-KTYB]#A.U19TI4 
@:E@5]Q94,3%-GCQYL4RPV2B@[#MRC>@S/_Z.(SU82=\ 
@T1J?)O(R;9NX40DX;2MLR-^>Z6@JTDG"%MH^,6#$ERX 
@KF3P3"T<[<I#;+0 -QIS?XT*(A2KA74C':80:.?"M/  
@ +DY58?_BMA[N'Q4<+Q2,KZ3%R@5;3ZO0=S)I/\O.$H 
@I^$"+QC'D7KP!;,:'B'L;;BJFK$!V'J=Z-G]!_R(=H4 
@CS7M4!AC@XD6=O@D6 -$] C\"Q0?'^F4)M\SYR/UNM  
@H]J<<(=D_J YEH<95SA2E?$J'B[@01TVV!;@GSHFK(T 
@_<((,O 0/=9I8\;I3NFZS;VOBT^=;D#&-<OV#K@!L   
@^DWL:[J+V,3<6)JF@N3F[L$/*<F/&@%P:A:6\@*N-J\ 
@\!8,BZRCMW(5'QOUWNJ0@^1,.C<:4T^E/J8V?$Y!P-8 
@1O#_?VMXU/@#"4Q:(XL#]FIA0XV%]D=I3Q(GI' :=HD 
@+GTE%'R >FDZ8H--CQ#/S^"TFXZDYH37_N(]()Q;2O@ 
@;=J84NA34X!"].69I+\B*A^P=_/W;<V"@G?\&1NJOM@ 
@IY];_7\)&7\($ RL<KD"4=OC\^E $9%/>6&I7I(ZH%, 
@J?WR<']2F@/9#]!#G@2Q D_!#0F(!Z8#30I NU:-:?D 
@WTM.Y%H[?=VR*.CM$_XZS=>,^-0/IH+&K79@($IL+$< 
@(KBZ*<-V"#A:"FOKR,V&'+JS=,8!\E4\2HU?E?:.95, 
@ZAJ1H#Q3-FY15&M;D:4DA9D-MUO2=Z0//Z5@FZ]QCJP 
@/E 1U(@WZU<X?&VK9F5MJ.\FD=/&!@#BR11Z3L1^M3X 
@WX>Z':-%&#M%)]/>7VRRR*D7XIAVU)I6I_7O7,X,%&D 
@.03B?MY.FGE#(]\)_9_BEKNJV;3"**V-65- -8[$6)8 
@GI P^ZP29K-:)G?&X>OL\S1,U@R23+8%,!0S9+)E0#@ 
@8-.Q-N ?'=F#!<\.Y#Y=K7P*C\'"UP\\>^X#:7CQ[QP 
@^S;Z*<2/L>":Z%\<2YX4-=1H&4>JSE.]70.(,8SDC7( 
@2_EUZ9OSP%F+ $41(_;+2*<-L3C,8=<ND(,6?Q-LB.P 
@FAVBV!OQ:^-25:BQM!) +;KU'<30$82_B[RR0R7HGQ0 
@K+NS%;VR'"'Z*(SX?&@XC:*O^;;/MF(C"M%,E/J6\Q< 
@YD%-CU':,62QJT"GAT_M0XF;0TH%B[F-R\ !::4&GL4 
@5)OC8*2/<]]8Y1:.Z 6./](8."RBE>*9FV%H9E_H6], 
@=L=1,5X_@&Y!0U3*W0 "!//'^>[AUST<BO-GT8+7R0, 
@1\%"H\F_FW%9(0E)EFA2O^RA>0'H#'(::2Q#@HOU7R4 
@NHK3:O/N6D>0=O#M"D<@3!>O<TEA202)<^&AE5!WT>< 
@E-]*7UE?;\V(S<P.%IWX:HR[ "IGA .#'QG3.3D\:XP 
@^.UJ[ ?8'&_H#LU0D4R$U0QDIO#,G-I(L1HB-0$: XX 
@RL"Y7,JI)UH,*Q:G2TD@7V_:_$EO@1_=4$-G-?SA<@  
@WAH6C_)P#VB(9>4-BQQF56KO0&2R2/Q^.:B, DDG3Y4 
@8UYA^(AP^ #6-!??5&6ZX_>50(/MYE'OXDW<EXVU](X 
@ 3Z.30/'WIVQR8( 0??82^( 8TS',CH.3#7@1\J$OH, 
@#ECY._3+-+H?K[C%#;L^?D'%_ODF$PQ-Y*JQ8":=O^@ 
@4H&H__@&6>/E4SBJGA*:7)%8W(E?>5UBW:GBFT]4Z_@ 
@!EC0XC% ):)&TI\UY.FW:2D(]HQ-G^MF12TN=1V9RA, 
@#K\8?:?@[[RZ.\[%?S7!5FB&6B [E*0[6)=[.8P=Z'H 
@;WCQ_[K1;8Y0\,)Q8)AS$4=+AW,]XD.GG*&!MK=#E#0 
@4IVG^7DB% H,L]37(/6Q>8\ML>Q-EOM72#K'N'R<H\X 
@F5%JT8R_ WA4B6(96>CY-+*]!N<+*Y''9!1""Y?-D(H 
@6;D3OG9(X.+T#>WZ<#=IX1$B."1Y%X<U!);663).R^  
@,K5<Y;+3^L#SU[W6P@O 4OOLB>UX@Z2E_PXGT?XQ3K  
@Z4L$G^[^*3MS,L:$^;OC+/S(+@"6OK6JM*;#$->$.Q, 
@U7M3@^N_>IO:B"L"IL*.M?]$3(=/2 5\H0D!W[#=QT< 
@?3G]M&E@-+Z##?GI+\MGSC+V9XA89C@A[X);TVAYSS@ 
@F$V+W(4XF#<07*_]:D4R:<_G&QK A/"UYQ^!>;Q)G8, 
@VN)^4RUF,Q( C,DS]#:IW9YB0!I@^#:0\Q!'S46*J.L 
@=#K%!AB%SZ"/;F8VA*\3,3- +A?;M,DTT(5QUO9M\*D 
@3]NA(_P8C-7R[U-Y)48F%67Y%+A:)AQTI@;RHW!/7I4 
@"M/U9QD0K-!_6PAB Q"'',\^R(O(17Y]^1T965G)ZD@ 
@$2JROPRW]9)%J(;.^0@\1$"$@[4D +%-+3X]9U8(\8( 
@DI.LHR11E99QWJ"QCK$/3HK[JU9JW3EE0B,XY[IA$ZT 
@]OJC&=$]*;?B&.3[9(_W[ ^D%0D$1B/8V4K=XZIT3&H 
@KZ\KDX)0VL7;V9FB_H(K;I4D),^YX,./9  P/5J$H,, 
@^D\C_@H.=@$QA*5[*:<13GQ\'D&Q@LPNBZ>6PZ6Q%/D 
@SGN_)WS&<@1? D<>!Z!M]AS/L]R"[T<H?_H023R%O\@ 
@?4X)])<O5>F%#@QZ^,7V7-CVZ!_%[LW;YLA72;8OHE  
@CM+[^;WSABZO4O[\K 5_D.$LP??)\>MHT> JP?ZF0!P 
@"U*7*6V0J9[^0;@MG-[_NUC#'?.(?P".XEWHE1CQX^D 
@<4M(,#V8H?"<S?L"FM:)TJAO5OU]PTO&8:,:@&! &2H 
@W E2T?^LQQ^9GX;@N'?)U98OXJ1VMQP7^ U=.S&B>U@ 
@3SI^.L5I*K:(?4[U3>V<H5J(.A8B]03!J/9=48&S^MX 
@N*7);5?%E0>?EM?V9/M'E85H%/=;Q\/;HV^6LB_O9FX 
@I(4T6/:9/,ER,<UA@O5:#_X/>$R))C>Q4OM;L<:1,Q, 
@;<8>,Q(]]Z\!6U=\>\@;_X/]\A,V ^$/F85\=$?LEQ\ 
@P[V5/+1F$8S][L.P29_OU?-=Y:"3+X+4'N)$*-J(0;L 
@29Z(IYQYEW3RN4>Y-/;#C,'./W:@S]H8;&7GN*+DWX$ 
@3JWZ3K_ZN!,9;N46P$!N3^"R<$).^/O_T"<XEV_S(-T 
@AYRO!:$&J53&0>2B]8WH!&)?CN<C4#\.QY,I5(_I=04 
@([O5W*H2W7F*;PV7HH2Z\7  "!)H/,*HP/F\'[K^HYT 
@I%KK'_;_++FXKC@:G9R8$%4UQ%W;?F%\_HY:MMG/*+D 
0<6)OW4SQ4Y6EO*>WF/)56@  
`pragma protect end_protected
