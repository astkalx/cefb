// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
knvAurowpKBJzHihNmqFzTKr6lctNASjsAJXf2VuROiXaxYSkmyGcg1THC0l3BDgopuNO/+X+lFu
WMdVfEWLoq/+HJ/IUegjKH1lxegsxj563Pqq4Xc6Vt5g83/1LPBfUi4W9Z3A24n/iT/2MKeshQNx
QiiDieqVPINunTI0lT5Am5cQHg3bOmlgSZ0DYrvMQlz82B6K+5UJE44vSFIbdEG569f8G6LTqlBX
3gtop6Ux5kipvU4Rnn7g/DrX6REjl9WMzEr+BabDBUxNPL0BIjAI2SRvY/AekdPlFaTyx6Xume3W
iBs1m1kHPh1Vy7fD5N8qH0uV2G97dOxqYThO9g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5104)
Z2WS3LzNEHYJG/FWQeqsuHZ4AKWWCQBq4/sD/va95JQseHmakl5eKdn10OV+wfK/1LxNGQmP5m8E
AYsnT4uL9FfSx97UqGa6BDC0DhfXGHEQaa3UcBcXmnUPnROYej0ggQtw3Fs51ZiBhBnwxQgPMVGw
IZweUbPyyag2XM0dh554cDvfzivhjsSk1m2AU/bn0E1WMDd7nB7duskH8V7ZzaxcKuRHWnXODirb
qB+/XDCifW7/NVlgMbdkOk20/Uwz8uml64LvaorjiZG1m389n1zSeGAMARDHWLmNwe0uHPTv68fu
H4lOCBE9ayAl+68RRbOexgxe/k6eNLMsqoMPaU607d/+1mgOmqyEE707rwnn0OuK92KAuh4LAs+0
Qpyu0HmBv2ohZBCwSiA8hvrQXCiNXSwUl5rEpoFISNq77pCtHTwn+EvsiVhxsrVn0CHx/Etk1BsN
gwPWNFjsDfbgy1RrBOsd0Z87Wlq1Vy/5pzwi4vsHo06vlgmJaslY1XNz70EBq9HE446uLYgOR4yD
e59YN1XrMNYXNb1/aG+V5LMic6ndw901IUuJSlL0BUdQxWA31rg6G0jr1OjdP3RPMRqH0A6z1bAF
Ez4MVeajLMrCZ6YpaX/OO7lcyQoWINpXTLe0Xvgzz9NxMnIxGiMwg9nrd3zh3Rnr1bgBxRzrmn5b
znNaBpY/8qe7cLZJzpzzVzHMAdWQ5lu1NW+TsyP2tM1DwEG7bGW3MqzLucAgsA9WcOIFXUkMHgzJ
d5cNwdw+FYMsNOgkFoUdRSQkstt8+rhOEgRnnNVQ/mHKHRWYar9DDc/uYU4+MO5YUv7Ahu1AaGD6
LhKHXWNpieCTjUGRxmCxR3xpnG8zmJPDA87zvL0bDyzs8WKyGzsQ54+MGTGhU8z+gGkFybzlyb28
WhNjU+h4aumB13Rcq7d45IMv9SOtBKzLNARu4r3bdYrIogUatwB2ollxzJG/TpyXw6+yZ38CdsKN
+h//VdTttCGZJseIRx4sqjKjA5a9s8IdvJPtuuByslZGb2czufBmv2xPf77NUN78hNup+nomS+/r
zzBQ1Qd9Sh9kGSdilmVdHgPfnqCd1ghGrxdY7DVLp50+RPeunpziI/vauiQyJUJgx/3rEMUtLbjp
m6vYm4wNWTwzyyXjYG4BREiTR+zKRpt+NSxbjSwAxoQpepnDdoX4rBI4/vbkrwJGKsMh34y9nuun
6TG4fUxuf/bw7XON1wEN+V/AHq4+hTerkfAUyo+hQQYAX4vtOY3t0AOdof9c26XigSnot9Rt3nyP
VPRXplbqe4z3f+sTffBUbUzO06g2/nT9/pHGw8rCg3SHlN9I8k7WuX+wik00JFxnkplV/fWLt5Yg
Po5VOX/sC7fgdEtH1qrEMWTb9jCMIf19W7fLXuA3CHRvQXLBMCuzBFu8Cdhrpbnjwd6Z9BNtDloB
DfYB9vBmnlmBbTqXsflurMfiHX0VDEBGoBXqWKAJ2flnRYATL97BVv9k56hUxdmuzwE4qFQJsYQP
tw1nQa2+etREo2tr1Vn9XZHTDz4+1bXceqS1IPlcHFw+vfvVPzgEOoMzp81VpOXbCs7Y2GbX8Dj5
igaNwehjaDDi9v9Qku7symTTOaIJu3JLN94LVu6bxk2rNfphPt1eTLxmblBuEl+0zMqVDO9//hpp
9Wf7I+BByXQoKx2xlKAyyu8IDFnrOmsKG+APj1XYsCfVX+9CLCEPcAjlG8ColYmivxAvgNY1Uy67
mO7YSkyDgbrk0RXmwOWhZcsxpkGvttF1Saqg/MGokGRAdcnwntES65Dp0RCcti+uS9kKeLf4kpOd
QUqo1+vFn2pd9w6IufDd82IwNmafW47E/WsJecrsssDJqkr3WUcUH7U+P/kI1uwseuapDR/15xa2
RpB4kGX8lVAgHrpSV8hMJzWyHN+cCodGMTX3kzvPN7p6hNpCD3GjTxCxkgPr/v9QOB6bPXE73lUq
o0ZQ+oUsVe8J/nQBEivhXZRlM0SUZ2kN4thkZdXcCFxORF61mdxXFKWZb+G/G7vlxVZqBcaA0PQx
xgr14atXSgn+qB4rdaHqgWDL2e4hWBLZFfg/hPDjR0eHwdhXVhdjRJUzB9NTaqjDehwemBJMKktm
QA+xsQEZTAgsvF2X3uD2fdZQ872d5PjrodOhyzaw/tKKOK8SQBWejyHyKYNKUOc7f86CjBqSkJTp
NZ2JKoDDTnwKEQM+IskykWNLkQEJS44UH4K5yx71tU2bJnJxgYTcJaQ2CE50XAVo04m1qYnfTUEY
KkXu9qDEO6WkrbfUdtKKsrIr7uV2TbTbN+DcW/dyHDn+daWcZ2uPqOlachpXyjD8Rutl8ZOfv0+0
l5v/CRSiwof9yJ/jD8d4esnMuXcUObajIZ8422t3kf5Xq05qPGs7gR+Hjgrc+q3lLYuCpxZKhhtc
yON1XGqdAOmadCquB1muaZbkFQiiJ91LPrNFFCuD1d4Rap983kTwg6fReWC3DHdUoACxXM3Btapi
A+QNEqYG+eAR+AnonMPStcYD8lCFgI4jGJ6PiUN5OOeMMEcXnSxIylBvYsuB8GC9rBWDicJyCwOw
eN44oLVVYh2d6wJbDNLa43zw5F8saRJEpMyr7+x4ggRKB6ShZEICYx9Yu0pR/FHbBaDbI1ZlYBVs
3PNriwGk3TlXQ7swc3gqCtNpSOFbTqdC4l+3RRQMHp+4kN2n1NBxq7u5OHJWLPbwXOutBOlBGxBZ
NcbJ9icVORdErUJG3zBujMeoNXBfPiuexrRVIbdrogCxIoSHUaZEYqZ+neupQir0kgdbkwL9RM79
zAPwl9P3E4BVSco5WN4svdAZ3Boke95KoEc9WkpOhUPhbdJauazXeLMA+YM1b8Ig6wqlgstCnqh9
n5O8v8xO80JHDuMFY9tiw0XFwFKKPtRI+W9ok0ISplTWpy8AN1tiyjxVNrk4I4GFZ8eermOCAFMZ
3Oo/028HoFWAb2EwGvTePhCmOfcaEgQthb84Ep+9MrxtGR1TvM2IjnCls+OBdqLU791AvoDd1SAy
TTkb02amXdD01cW+f9wnFBA1PWz4Y9yNArOjQ01X2wrlWwUGDic7466C3KG6Fo2n4qbf9VQIMvyc
LrP5dAeFONTt9/VQkoPg3GI6iZ8q9JFW7A31i3EMoJsW7ylpCZULdSaDLDYShmuOOLWoaombJGhh
sWAuLU45lG0GfUYwtRC5A3sYo39y5Wf3scbtFzKSgI9NBpMttbdZJD0NLcnfmxAZcJz5ncjJXnGC
MYugR2A21KtPtKNd1IjOLBJR+F/2KnKfMW7SujYh+SoUcl32BxRkQuWeR6YEPhpaSJKk2BIjFAZG
7fLEoiuhcG1dW/ZIUaGObS5o5ec61dM10hCASnxKYICcwB1t0XdSGgZuhg9vNAWKMeLGBVWz6LRl
kV6TPrrxNb5pVKv658L73nInylIGyxzLZExcu/Eg0BWvL6PuMk2A0jRZz7Ap9dCfWdVuIlmp7hUa
tk1sIpsqUuhyLEPFATHMDxftDJ/XZfEU+6AzqX67iMEkdvOqjWkPE2E44WQ/Pe+VoKNlStG99vDx
4AG8fx/SZJNAGIjrrn7eiFcIxFyW3D9SXnWxP5HsNIBFYkEqVpZGI+chuCbqamEmGdGZIKkuPEhx
/x65rAbhF+aa0SI5ytW3SDQbUjElb0A3RANfU2rEn0m6OMBVBxGF78/YvO/e6ByiOmSI0xtCq4rf
ActhQ/oAyRIJan7p2bzXkUXf0uk8C18aJ1CusIfAywYJhV1jbPOfOxdqoxYJswlARBfhOhrdXPPa
uQt3129yYVqYRgscD0owxWxthbrYqdvGcYZpmvClaTr9ACO5biYht/uKTVfhedcR67cjsuLCUKYw
OsNkZkAO3vTQq0DmXxmr4OtupZuEtn6FN8BOLNiuwHTAnd5amVuXrQe0gtDzVhBjS8EYVZtVXZPA
cJyzzqkSj20uQJMubAUS6HZx6JjM+RR3Nc2auODwKz2Wp5MsLpsb8AIQLtJUVTMBInhJBvXYPUyD
dYuRSvcOO1dfC3qpBxj3M2GfK8nD0qLMfvXeDtKnyC9opA1FnudX+Ga6uA2G/BeUIAgiA47csB3g
TuzqC5V/UsTQjH54BGrm92QUiVfehg3jdRyL6BxJ4ka139wxF8QHQj5/ZaUSjmPIV1tEPIiaJALi
xf/GFymuBXt8nXde+d26d+At2kYDXee+AqCk0ytVD6sf1pStMj+o0IuL00ECS2kTIfxni+6tyRwD
wmmGzHFM0RUGSbth4jDEBMeTsxTQ4u20uky7svZig/+MbAhXknxM8z7hUGT9iXRnZGgCtSsYU7Vf
eCkI2WhBQn83PMb6k8VB4QJUHrmF3hZlfCTAkQYUX4ZCCPPQi+WeEihvUVlkftCQrA2ODHg4l3od
EzScOcJwNszErb/oREX2Hh/ExxuQz2SY9nvT/tTR7zNdFnHIJCrNzBXS4YzFCJ7Mw/cFX96+OYGo
yx2nnmnSCFbqFU85PwWpjgWcH2ORcPiUwwHv6dKXDv/AiF+NGwI2MwD3o5L8SPb2hIqNRCkWNiSG
QQYuhCoyXkvQ9aEGt/Qws8hUZnb+5i8wjSVk8r3N1eIdl5xK511AJ33GCi5o52YSj2n4uUepMAC1
WzQDm/nNbXRcHUEDcP8SmSFPkZzmZTRWE77MxbYYNdRgDWqg+VwV70OQsRy8DdD367bZ72llL7nL
DNj8lxzcX/58OkuNOoulLKTL2ymmCJN2TpimYFXDsYd7iK7kbY5nF090zqsVzjt1uKVZuh+wdqn5
2fiCW5c/u86pRz3H9GLuLw541vAFj9qpBhIu9ZSaJG9bU9EgrIBz40kwW+/tlS7Xcv8vEUk4Wcjo
7oY3iZDPvh0XozpJ7VSz3QNv3AL/JhHFN1Cow2RFLGvD/JMEShm7mBvuwEwGyQ032GaQVrewuUVS
UgAzpjjRONa5jt679RIqTTe11lv/hH9WM7isKB8vV0mraCPNEhD1jHYRFTDM0Om53bG6hVLoX8QC
AiJ0raC7MJDROUuaOjYjlzaTQU+wQ8oxo8sUOK9HYWKNWDWKwNsBGMZ9uNMGEsnzBlW/YSKYAq7h
L2X5hczgboovQ/BYqZoczPqWtGJAW5OJFgt6612312D9zmxF6NL8oEw9dNjoV+uWfcZce2eDf9dD
luRzxpPVWtHDlyrGsLhwfu6MiuM7YmzwgK99j0LaNBodoCOO9e/ULY+v+B78q9FMrNvMZyeMz1FU
cxoHFS4w1bEQuErjHYw+eGcJoL631Yoc6exVarzkEH3hNuVFZ6//UCOuQTX912LZ+irGnVTFqhPL
AkdpND8jzBXnmYwrjQMpy+JmmEwsG9ENpTOlfCy/1kX9vDEbPqXakl0QejILohbQjhDo9RnNRrb+
mBkT2hOtnoT+r22G4blsY2V//Fd1ERU8ybnyr5nVG/ohqtboPcoxqeK6fRpivrpz+ctv8STaGvBM
OkqOIHTdnAYu+WcNDshYKBg/Sdo01jIDd4F2D+z5XkLlZ1s6uegMIxOMKOKW9UMtp6vxs8B+nbi4
zcIo+45LCPho9wNJuyRGgVmH+egTGanW64ng7RE8WlUgTVzynvBzdGmv3kyQ3mQdoUkDnUnl1mIU
H/MD6V+s8Ong+YcY9bxFMCMdT2azFodPdvdsfn0zS4Kg78lhOVzDsddQsuTEAzD8OEuOHEDirq6J
su2Y3/AqzaH4+ygMVnIuARMRFHjYLRXnpQyzmmT8yCoUCPPvdoCSdl3y73zneXnwZEDnaN4s6rWP
9gJu8bBdg04aMTTUUFjh876a3ol+UwX8cFOseGFs0hA/8uhwibcE04gLibuUSUiJlIzOT0He3OrD
I5GXgbIFgPSQucj6OtLHCXs1CkWUJT8rr4nqQPdncihvs5mALjC+De/iZ3eUUGJ4xdyTAjTWy5Kx
mM6dTvr8pdG7PNeEuMYYwdx8znhQkdwJXCLR4XFa0G7e799ksU8VPJE13+5VLEzKqMhOtLsRcpWZ
SkkOWxW2pXoz9KyiY4Z/fkHxfTW4yvOaNmS5esAkM3qphQxPJnNeGYMvpouuyM9tbRLCufZ7pDhY
MQAlecIErvaxmwG4i4PNxraKYO429RdUJ4g7V5mQlNs/9wZxmh8DYp1TV2OH8oCm3BATq/EMrxEz
YhFHo2IaUa5KpdtsbWzo25N1aKhHBsU4q6prgiuMR9UiYt/AJdBSkcOdL2oyeCwH9lC8qWFaB7dU
NCEBawADPnufehK8/mvM4FZDCaPqVsn5LeYlCwF8tU8MYecm5cvpB4Sh9tYM7f1dV42YkzS8cHwF
4VF5GzA6RyzOee41OUNM6GeYjdu42+VC/5AFbLOYTBBOCCh2wR68H8il3a0BA9g8xFbheXj3p2FA
0YhS1IkDZ3gLSN29zIr8205O85ol3qBZS5GDQvEpKK5I+gHXmoh88RCfoX9EnFKZzaLziI1KliBd
Q0Ff9QzkRBoKZVVYvPiBi5yqZDpGNcHFMbap4MwNR2whSo6Av/RBpz+QTU7w6YOVCUjr2qrYLffv
vF5uDo3HZaWnSPDjbquXkcdO1U2UPsmYn3ch6P/+NsDNTsXd67/Tr5hWjcZzqc6t6nO12u55EymI
AVk9bZ5Da0+jcvUmoPJ1xMd/6fh5nLs68qR6auU63UgcPl49iBVbjrsKXB5fCvwYZeIAsAT+ARJD
M3qaKWgYFfOGwl41WJYooNMxGMgejccH8HX79Vi8ElQV0F8XwvVGohrPfpNwJckNMVZAa3X4C0Jm
HzxFp0b4CleLoZSl9sz9zcYsMlqN2e2LTOuI33Oqrg==
`pragma protect end_protected
