// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
nujgYmNztCBFuZQTCC7xoLEEjJE7s2eQwVuC5x2or1mmCIhSiyrji3eiHrsXWFdZ9J0owSuNY2MY
vXwz2U6w+FKipKBA5tH4qlNS+ztAqInasTWyQcoZfguQtlRojsdhAnjv1rrX5fVbJe5v1zK/enJU
QIZ3Zvl8wCUAA+kOI8rWqunLHOYF1YoaP0fCdFBokabL3LgAtN1TzoIo7NoBUE8UikzBTF7KhTe3
dqJYGmVWVLrwtWwmrBjdGxKTsO0mctYB19zeLf993gdpogaRdu24LiTkzhYjYTf6wde5RhyYI7Y2
JpTIMnUcwjw+yUzCUou4X0cMaIQzaTqju6ZK8g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5600)
BAOLR6JxrcRQ65qbusrdS/JrcIec8qhVPVJIvWeSqid+vZhBfx8YUfWIM+4sjW0uAo+romX/31uG
H2xuWkYkd7Io7SiToscr681F2b2q53iGTcA0bwOYIGzIqytBuytbZdFYM+pnnP4Jmy9l+sifHhR9
u2ZTp/ZjpEoQjVOy79G/GixEq+AEVY2MCOU8Hct6csAOHGpnSNuF/TzZU6s/Wi+Km3pPnBSP6R+y
UdUpYmiAmCQ+oa1pEnAgqxBPjQ6o7pCjdtpsRaDVJ38OZtzTGldKkRoAMGSd6Vw6W89MIX3m3J+T
sYLg1foch+oYLcWsH+kiwotW0luiUQx8eHj97SDaJFip+u0IMdX8P79BaScTKAOjtYLmIdDMCJCD
8d2SgtSpNziZtmPeHXtQ1Uh+6EWI/R4/vNV8im2MKLfwueRy62vt7QfZ+wmJ/IDBmv4gGspnkLLh
ID1WfMAgVHLDdssNi7+yxDZHcxqoqt7NwnZ6jpxPIVmbIbc3gx5BbF1bObFi0WY4tSEHLHD8l+Fd
sJrNX5Wrzh8bgZRHWCYQyIjoM80YZGzMohCtDjRr8cOzYPaqp3+CpZBHBqPFnHlvUpUxNGP30RvN
kTMj8cCul9/9024SkgwTkV1hKNCbCkrlH5M+cDHQFbrOu06oU/Oxn0m7qjT17FqhKVuIA8R6JlWX
ZJVEzK+78ZS78QeuS3W7R4o3FdM9mPW22feKMukgFpAo8phdFI1+W9OySD45kIrU3QgrE2DCHOTe
i2CATu07UxNEU8NhBkDcqWVkbOE4yRmlDo49JQ+QZG9tC32f/90bCx2Erpwuypg4Lgf7bZ0PkMAT
BYDeb2LM2HbCplvbmXtAp/LmbV4E1g1TJLwNfXExG8H4nmti9qaH3qom5290cmhIO36LyZkdhxBL
6eX/VikN4u5oh5rhpVOxa1fmAASdJpW52A5B9fjZEV+DKrVDiuJ6CkklCY6DdrZIlgL8KAjoPgRg
IaRhDKLCPd4cm8yfU4cThJzRu4gCqQMqCaXYJ3zjaGqaQfDNy0AwYmRw3RYGoDqQ3wkvb2njFwnq
W/CKtCbEa1HmlZHXM82SSGa1KcVhgbACLlhWM78GQUNY4iIRO5wHz8dQBOPFaESsxucOogTxxnX9
xIu5Dk5zDIAXlLVAN+U3lkQqjVViM+1l1RNj0Age0P9h8v6Z29qwyGVx91sYV9YTfC5kEOBQ/IIg
BAllJUr6BQzxvVjnc9dyfYsxSlBCfW5enqwyHAia4HYudROO3NVr6D15/aETqWf79GbL8xc8pD9j
I/iSHzs1SmCi+8Dquof9kGvI/WFxTQ/hoRxCkaiTRrBREWELosoOuNmf1Ww1c9IrYGoGaLW+Zd5N
ETtmWKLEBRtSSiTcdcTwOJd9lWrkxRh2pJQLsbRyFGBllBPkwBDT+eV7Mg7TfsrbEMEyQl5nXq96
38svxOQIoJSed1MQeKoibyWSo8CsaKyr4YCY8FV0D5JToPWZkiW8YUwPdIup8cKbhYNhf0FGT3ba
W1os/bT25a+KeyZTB1rwJA2ADNZem50wsPRR+V6FOaTKZB02sC0qv5CVe2HbSf1APrPDLKUa5uAd
mFIWG12O0VytifgPPGue+9+aFa5WUiqV/kg6ImtisOhfaAUSHWgpUjsC9ZIC5IzhSY3EdMVDBkXJ
En3JbtkEmj1GocRNNQ3FHO/F/qnk+Gj3piYn96ReXVAvP3pgZoCLXdKDFKQmtXpXBo5cfgfLM0Sn
F/e8Ch+SI42PiBBEE/mnej7+fOp6cOduaJvqu6uXYDqw6RN6wha4KMKuLUl5DljyLisSogzC4Jpy
Ny77iwI6E9bhN+UqHXDHFy59n4jzOeTTwbqmfA6B9QWgGtdBRgec7J9CeLW7xAGq5E1GJsJ1vUTs
cmUI4PdGHQFvGs9B0eD4bU/HcR0ggSh5tBfrHZC9qLmeNowSF0SUp3Ru2nzYoltwTL6BdAaANB6J
eDnGIRf430z8b0UiU5+aaFZqMo1aKJs4c+oLAmpuhxt94MBcBwnY4ZU5dAfIUTvEZ2vn0DulltbD
YNEymocHxwn+Qq3ietG906uv66PLEisO1i2Y1qbH4Fz7xV9dknTaK6tNukiDZxTNiK7GUECYWiR9
ohdhgQrJdf5zFNW0zgfp5nLSRtd4TgQxhnXiVyvui0bzC/B+u5CgBILsckSS0ZrYz8tjFwlEvqcF
R5d7cVZYLWOrUDdh/8k3q8LK6LztuHMLlrs/fgtEQQTLbtbycRDo0zM6buAlfG2HsJIgu6aSXr65
aHEju9SsGrr+qzVCJdjsaaSvwUqKLnhVwPZgPZjR4+nddUtU8O5k6PjsoQ5E5dKxqEj03J5HCk4h
XoxDXEQefaXawA89UjkaXiKofEUfQBwGWKD2vhGVvavJJKF/i/Ub7ABFnFLhUrJFsyvx+C4UIE7S
VZpOu13FKwsLD7Fw88y25SpiikHlNdrCmdbX+84fIkV95SLkOcK/SkCRHqoOp50Cgncn4NCF1vh3
3+BJdH8p0M651D4O5+78ITFDerTy6xdCIIBTn0hRbm5bOZY2B19UA2XXU1QXvQ4IHiOdKmaN2rem
63Fi8qkQO1nTRyxSKs0JzFlBq+BJyVYRSFsJVVC9kCyf4XxwZTTCm1KDzS6bXmr9h4gkc4YsKif9
bPrTsNlFboG37DeQZPx4b1HRO7MtB3mDYsvQhp53LEvI/SGT/U6ny2kF9wB6N5VYzrKvBeDoOfa5
aEwN41O7O0lsWLPqZi6KLwgaIYnYrmJuqFTkvs3lS1z0xPOdJG7aQSZlnCC3G1O8wFemdP2rEIzH
8YK8K+PalaoCnWA2g7Q6AF8SwfPx5/jk1IJwSqJHKVbVpshSddk2xiprNTkIeXFH2v/PBK6xjp0x
gYV9Yp1BN8WaakbfP+byv14bFgV2xx7ne4l81+liOjFMr3xuWVWsbOyDu/VL0DqtDwqqiDqoTIuA
0DaR9Qmo2MEFMclclYgrBjeHVb54ViHL7BSnwiw8rf3fgbeNAj4a6qzDTI7hBsQyzvsQChYUdSJp
e4R3zOMvY5d39zXpSD6tuR74BRDB6gE7Wb3/LVwqf36SIk/yBwuKQoXOoj7vdGS5SV1PO+ru5w3m
pU303eniMOg2N0MJ9JRIhgej97dP+B1tlKIB710JM8YZfn7ox/qH4Ufp5qTjwaUHwK2KP5iRdkhE
kDdkkEJvtNNi+B+EWuVr0cCB7wmkOUE4ejYtPxpA1wG8G6DuKHLdDJh5YiepV+3HtCgl/sKR3VlP
L/y8/di3wHW4jEroHA9oms2xmNOc5lfTQExVQyEwA5PKBxOB1+Z2cxrpHkAlzrl3Xm/1k03kEUpi
Y0j0b8m1G2QWdRxN8oFrlZYWBF01z8ha3jNTtIneE9Sc6aY+qejET41XaF1EU22A2/Z5z8zBHWuv
IKnFp3+LVG5fQiJ0ZKYXyLoEPIZcpxSxzZZBGmbsf1AWr//yl+sG09ZY/0gyDy4xFqqgNnfWUcu0
zIg+50KveacFz33kuMi+N09YVkt6j9ueddrQwTUgj4QzOz95oW2jBhCqUfpDV5hEW/aW2QwZxrhx
MHjPX2Wd2JklqpmjC4hhBdrY6y4COQX+B/baAsyjbWG6pQ9cA8Xf2AUf/HivQb19Mfqt8jNDefNF
4ADOUjOgyqavyx3VzL00yBZHwZGj4cpFRahpG8EYNkZ1AOckjnGr2Q0buM7+At3fqyckPqgbZdg+
4XOsOnXlfWnVUb6+nfKpI5lE3i6ecEofnyvsbzbssTWGSpIQet/kLFS4y4EcrqZlAk6NX/jaYKML
ZR37Nj2DbqbpBX3iwI4P5xPZyuuC/mpzuDdQyawqdmful9a+wLlCYjTtD7Bd/8JvNULSD3XNo4uY
Ywj7tzx+RC4cZMK4D6D4SUOA9E398gpqO5vWCUso8uHd4wqtdVnF6/Kp5O2zgoStxfhcMUQ8dm/C
7g3lMg2Bx+bv7A9oaHD5WKzP05//VuqBQbL3+zaAkICo4L8UNgZCXocXHxaSHGkE2bQflLHH+Yf8
KCqC6Ao3fZXuFNjoDH6R1xfUNycb6GGQzmukqeSCQO1Lss+e8BQpNy6QczAUhmTUseeloU+AJvdy
KxMEjDMJKshUjZuKvY9HuMwOeL6KGwbPUegFSJ+qc8qN8j7M/kOM5x5PvfwD7KDRybW05pGBhSQY
PSPgREpweYN0/3wZllGDl6nmO/9jOzRrFp3EcXIeq5Ms5zq6bF5vMOqlwyEfTWMRyh1xj1mKZUNW
Du0yOOyF6U1xpNlbouL4z0XNDUHa6yH9N5YPLD3XTrIh8OmMuoSPDgZswJTlFkfhrJuUvNS9kVBV
q9wmTIYyWJTbydUMEY+dEGqN3xDmn0Vty5Ai/Wp2tuAbwNsWufwPpxUjSmhWKm7q/g2wKSlOi7Qu
8OHeH5ez7/A0PKUevFYVjOmJNi+XBou34mAl5DRyggi66zAChKE8JSGF13PM75e887q0EyNi9qs5
/9jEZ2ZLcKOFWwDNt+iFJbo/YiVH8sl6oFSDM3Mlyay4+pk3LkUpuVQTr+nYgrzaj6shVfCfjGdb
KiyuztgsV6rlvICERYrLhAcXF40CoZ0151Ym21Z+ctvmcuFr64fnJcDo3ybd8J1/xVj+uOxS6Lze
1MLB1BjsICgHCTNrmUC9HYAG9gYpzttUtlBpjHolzHlS/atG4U4ZTjxXOTCHSW4xhlURG+IScQUO
ASUFD8sHtcw9426fqYjCtavPYkV0RAMQndLVZ9XfnL2Eb+uSNMUq+SttdqfGuTI/hAKpGveShaAP
2+JUwp6sC/dEvxYNgvwJgkgEmIsdPYu3xGnz3JOV2o+ZrXURXl0gmtBdapvSmuu/XZrSRSYlBRwV
XzWCRsjxt2tZ6W21GIldQ8gtxO0UgMd6bxsmoSZgq7TAn7kNPChrCletYguOLfr65fsXWKx7abY/
CAbEJN6tWbVyx/aWKHy36Uom2sCAY0Hnw+oms1KLNPnKL22YdFp9z9vH4JF7XqQ2ouHTaCoMCVoM
Nn7z/zI6AENboYBVHKhgZ3EP8sloGe6wwnrWMNimIpqM1l3Rea7OYUlC+16jC1M7Ry/ibCum1uVt
K6ujdnF4ozzHsptHuKRh+Zi3W5CMnIPaVtU2BT6Y9dKEpFX90f/H3fHS1Ddk/f1yYumfZFbOm3JP
bw9fJ58TYAgVjzZ0PsJs3GOGWBmQmtfYWHcBGkvFSb/4dpafCi/ovCFff7kzOa7eXzxsHQWXjAaa
nTqJEwHBamH+6EtPBycr0XhDMxRgllHZCMll5lca9kvCytBq0iMewypp2Kf/8+bfSnVV72lnb753
rD0XGCL0Sl2PVpcXilCgGzU1w7FW3NAdZ28r73yJmOg8XkMMyuG1Vzcligb/LyZtaeDPxXjhyUAE
pbqsngak7o2h7LxT9ucuGIWfb5D+nt71ifgMm7aHHE091VxRXd/N+U+CabT1312COr6zx1RLW2FL
jni7+ZGR4FvtQsAwtksBJlq/ONKOY107tjmr5kkaRMp/ROelMT4xJd1AnaLzhPisRrE8oHNJR8Qe
69R+/Ub4SzBqUe0aUg7cXzXcOXryMLwhzFAMZhew/moznae6MyM6unBJ8X4avDoTNc4h4Ozda6Ls
dWEhVFjzUjsXwH/W1iJ5waNWLi49j63YomihOhFYH+moA0aAYuPhngi10PVE9c+D1IoGZhGRvm3W
ft2hWSJPATcvVJU35GF4r4sUomfdXtxmiCdMnCorK0E3/xj+etjAeXKyJgO9BR+5Zj3YY2HZAoYD
bkEPvruPaD6QeXo0iEJNYuzbKl94FN3JwqX2lSWIySgQmAD+GooDNSAKTW0YQzuI4+AE+eM1GTCH
X1GGVRoue90PpMozD44QTZ5yjv3BRzD/+/LA9J9f7RM/GIU2u/7DAGtcNB5X9fmAYT68tKCE5FgW
IfnqhCCidMAuSXDfqjqnUEWihzcHg8FSQQe/7qfQRkVE3TnrpvANcBD/YdrOM4WVmbjDJTAoPw+S
yY1PwHQEyeIZQNgnKdQEIIobjIoZ9vmDqZ1/j35DCLHIEjEPEFPT0lThKfbpT2oF5MuoPEjqkHmo
dTjPC8OGkgD1vO72HpPvDZPCuDk36aqmK0/1pI/Yr5FzezQn2PIF/+V4S6VhPQ/3WbpvVQOEQBwY
ac6OPaooboIe9yZbl17pBlL9bDPl4WOZGFjod03UOjT29jW+Qej82O6OYCqixHKsWxkJ7kybX4af
2yHVVQi1vhNF7x600KF03BWs1qUvLJPLTb0FCmc6x6bHMFgk7tTpSY1/LOihUqAU/JNjX2vHyYlr
Zz6ehcWz1cSuhe3c7ZkzTeto06r77QPzO0FrgczIeEkrUDPANLYNwqNS/zSswCVeu9Xv7tISijsY
kYkaUgNcdgszzhK0fU26lUV95NlEQ387TeWHGbxrpaGFerEBL+Q1bPVo27nslHY9G7mhM88+XH0l
msrD1WClnm7iQb8D5i+umJ/YNax7YrgK0ZJpET0+MdpXutdDEmYK5RwcS9i3cL7ssUfNqLBZSAuj
TrjbtveYYJKziJ11fw2MYY85NFP/Gl+HexlAOyOn6f7JJKtePV4PKY1G1O3A3M/OgCigOOfalhmx
Z/p7TelSZa67dSJSPiLc0CCOBP7yA6ct6RWAbL506TP7xrNNEOHcid2V6EwQRjbKsQiiwjkuZV3Q
h74CTsSCAkt+v2XoVApCvTwrxGji37rzotwboJVWS5TKtQwvg9XeSGclP58bc29Zjzt84LX33GJr
9+X3sjpui4obrmOIOaLUxIJqKg2FxqR6SgeoaPTsuztD/30gCiRgDsP+dZPbw0Y0MOcMa3CYnO4Y
/pbzFq82w+tUiP95IPWSkT23ho5TSBHe0wR97Ad9eEVW30TMq31k0+umzfpS1DbIwTZeopXmlcfL
TA9OdaeInNH57oZNAikVYyE4neRV7P6JqIl0o5MO+FfNH+c2EAH856PbDCuoIYuvQ28Iw4wp03Ld
D+7Lb3KIDW2bRXcJJeMBwkvJbPK21yEpq+GlCkJhWun6B1Xa52RLzciHjRwoGPEkHlsFHmrIbhvb
6EVu7QS12hKEcBqacBcMgumOQO3KWMFbAIpKsTlA/4agZsawt0sN1fHTkSNLyq7Xfhsm/T2V09wZ
95b0hv222UzL82sW5vsjIxXcZQh6yB4TGquvlVlMcCPfQEQRmUMp1VOFLMVg5Z5f9JcATbxii28m
WskPNwnGBG00YqboqiwbIrXHMZ77o9g0etMe4Iv1vI5Vndulr5RVH2EJfpCVXt749x6GMnn7GE3/
HqjM9le4OVwRgwUI0tkhlziGdJAcdW8kMi561es/aio3aP0IZII9f96GF3IsBVqLpnarJiIZh9pq
Z40/+NwJ4DJvcQ3C6sIuwVOUlsmt4qIwNAA6hQgJoqfOoxbHBs6kPpO4gRJMnm29vcGlw6Wk/edo
Iy+e+a5ZPzXknaTRoTY=
`pragma protect end_protected
