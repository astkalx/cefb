// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
H._= L,7 SB5W>4EAN?3*C^P)L?F95D.L]C&C<":_C>ZXAOXT)S1,#@  
HJQ0-YXT8_,P3?ER$?&L!7J9)S!_)TBWEZ>5="=S2N@NVP"E8[Y=-1   
HG[L&T:)NM/Y.ZHA$Z9/YO?<*OGJ>W\K;D@Z!X>Q]7L]T'9L>+2O[^0  
HQ\H8TF-I41B^L'C,&N "/'38$\HE+(:[9-#8:AV%!^P\#KQFZONM%@  
HKJK%!"?&-,<WFI<7W8(+(ZO^?8JLXJA53Z34#MJ^J4IT$'#3D<+WQP  
`pragma protect encoding=(enctype="uuencode",bytes=4464        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@=AU]P'H96 3U&G28?12 5KIZ;NTEW4P"M;FXLFO0DT$ 
@.V,) >$JD]T^M]L56(Y5\Y5B'*"K]\D'].4#'E94PD  
@/4>X8J;YX2M#6$8\1G^H5OG\ C(8'-HN4<7)_%M5%=T 
@M9*G'^K+8DPUXS +3*?C_<,1+,A7Y*M?@0V+#BDQZ\H 
@31/-[:6B5=K[>2/3KN%!2P+J*JK]*FJ%;DY>!<^GD=\ 
@[3)=GKPOG0#"D"'&WOS/UCF1L2BOK2YHAB1CU4W6G%< 
@?&C=)8O*G =A5*OV,44PX4FG:B\JT%N+&=*NL1;ZW_P 
@X.XKNR$$L=NG,3?]#+-'473GPJD-HJ%< 3V665:D1:\ 
@T%PM01 ]8-Q:\848SN]+2)&+B9^\;"U[1Z<J9J_ZH^P 
@^9=G:)O:'SR298OQ"JC*41424WX6OZ=OF&IONC7_1KD 
@R5UO"%/DLLGBP1<J9*W6Y5*(:#$M-@7TJKN26/W!9W( 
@2FHG'/?XQ[N3_65N(;AQ'@;-G]G577P37;CN2C=:#Q@ 
@G]U AL*"'FCSJ'.'2="H_D80V[ND 5Y#5$!5-W^IFM4 
@[H>3'GYWS!2\OOE%GYSIT8J\Y[T3BU\V$X,.V+27OK\ 
@.<T5<-F?FN+&8E ')WTJ+0/+YO0^)?VIX$6._$ZZE6  
@X*C"2G_RRT6WEUO'&R[*<:YDL[A.DJ-+4WAHQC]'OD, 
@8J</?^IJ/Y1J+% *BUA%\ )2I_H@E7"U91=QXYSR0K  
@)V(/SA\/?]RH3&S$%%6WASR%YOFB;Z9+&KC=%Q#FA?P 
@%+T!-EX\L@[%].F/J\E$3(TF7D!UVH46-:9FW).;!:, 
@Y1L5W_^BW9LE!WW#C$C42Z9POA!&D2SK[RE-(=^@=K< 
@Z-WG 5+TP8:.*;T=H9'IT15SB4<E!(WF3#0A-4!XL>0 
@8]=J'XFF/(ATB]7T;+<]^8/0)L>M8213GF?*@L@X\2T 
@#(5/W=%]++=P+\"/!X)[4]+,A):M[V"\!;/F,>U;7T$ 
@9:6K&]F[@$\.'AL>$I7T8=BK5&7P(+UI0YM%VJMG95, 
@<818A[0L4B 6*)Z911 ,+[)B8C7T'<0"LP@O*3)6X>\ 
@#O66)5W9WA%54'W0.E9E>]C)=_LFT_JV+UP[I-,#QR( 
@0\BEP%PRR\5V4LZ+*.X8@ \8GR<^;W$V4YFM&#-;B(  
@J/H <]IB'C1T'_(>12R>;BJ71H\%')?H5K!]U_>+ <\ 
@?P<4XI3(3&B(R$B=ABG=U"T826M4/;CRO3?:H4O3I+P 
@DF45X-B[NU\BX!R?!$L5(!TY. 7EG#;+D'/2V_TKK=\ 
@1PH0$WMU]%GH/EYBVN^J _=!*F"SU=MR2\)1S.)-O?X 
@2%&($!1H$BSZQ[A=G,*[$L[B:.EK!3?J\IATW#:#$PD 
@+2?RQ/1WMQZ,E_2<Z'FSE&I$Z?R'$"^3O!5Z>A(-M(, 
@@WE]E-Y%O-N@F")U($Z0)CFR9LR&J'L8 >U$(:1;NT@ 
@O:R0.,/TTTA$=+67)$! \XK<YP0 )1;RLX>"O:\MG[, 
@O<7\.LBE@.7::#A4/_<_83EN75,A0:)^^O:/8TU;>B( 
@J0GKUB?-8?<#9/&JN_"D<CQ]6HFH<%O-1E\RJ6X+P_P 
@O9W@G3&0[UD8D0S/S^@B6?:N\7--@!F^)/=SX&\!6"D 
@$#E,=D*9)<#+.:"IW19<@AEP0^!6JRV$W8D7QI*97_( 
@4-5SKN='$LN&]Q"MXJ%M\3P61 0U")"K^QZ&Y.P7O24 
@?U"-I>5( O F)E2$ 0<OV5LX\[Q4.09[YG73(N+5H%$ 
@3 >&T '_>J9\!2HU,"MFR%;(HF_T;;PSG.^L(ADH<F\ 
@("2.-U7S!5M!#U[?85M7U#XD_L3%L5@?ZR==\"+"SHL 
@].W*R>V07V/NOO/4Q0.6_<'L/W6"/P-M^'H'8E.Z#A@ 
@<K(7;W]<8)"ZS3T^K_EDY9 &T KD=/BFZC;3-(-'9;@ 
@6+\>Y?>#[1?== $4[QH7<YBVKR*';3F5A_'J16$4P T 
@3[RE[R]U+*"?+^7P6]\ULQE=U/VD8B$(*VMV?D_X2R0 
@Y,/+[8\P.'$46Q-L9*X8FH4)4N,\<1!D7ZLW]G1G "\ 
@6X2P3LRD.&(2X84,-J(^C?JQB!Z[=BTOPI8G=,CMZ6X 
@JA#J "!^*",M&YB7C8=W(>A^#K.=JHR^56I!*V!>IY< 
@>4JEF02?Q%=!F=N^Z(1".HS*%Q%:!^M% \-0::P";FP 
@2U^9F*;UNAJZBF\U(ERU!(>G? "PO.ZH \Y/&[&N6%( 
@IAYZI&1'4,L_R!@RB03M?>_AGJ8CV._V0_F]^2!/Q&$ 
@Z]+5>SP_\%A>I/K;<D!S.L0>"I+L23[YMWL=%DAZ6OH 
@[P_*_NC^"63.T][Y.!O-UK2^X]"A,MK%3EA?W&<9TYL 
@U8\-<_",)+9?\K_OAO_&'2?;)=^SR RL9KQ#U;($JP@ 
@_] _"<'X\[QV( G2\2J7O_5P9N(TWX39' Z+/#-G<OP 
@+[S$3.M^#&'>^J.0J+!*;UUT?6(2 $H& 4S0S]:N"Y  
@^A/.9(>)Y>'?.1_,TJ[J9^7#M\,@T(P8LO0G= C8Y@4 
@=A]E#OC4#3)5WD]5"'93:/;Z>5>#7+LQ<9S?K_K&A., 
@FE32L@\Y^@>89>, B_J\^, 2D5(ICU1I)#45LAP@IW0 
@GX1&BWHGFN7C;84Y+S+$C0%[8;E[]J#(UNN<P"$?=Z@ 
@P%K*L9.88:A_$^^\WG=10$QUKG+",]XHL0+_/!!XX>$ 
@%1SJ WL^L&HV(_5^+YXD0ZEQDV#MMBUS$4\L=6"XH=H 
@<36&6"HC,=C=:!^_BZGO>XE<OW"S7K,-4\P@<IF@Z%  
@%:A)V\0+<[J7CT3VPF,/V*LKHT)&/GN<;Y!&Z2B);GT 
@7#53,,6/6E+I4W<1GI]J7>&"X'=]8@5M!(/ MR.+:&( 
@ 4F^O\!/%_FM$B\Q*8MF]-3W5Y)7@/][+5?\$F+'I$X 
@Q=]!S5%6=.>6YUZ^I34;.=R^@*EI+P3@3>AVI-VEDP\ 
@B_X!+*#+=N'%7^>B_]2H:F(62<*8FW>:9.;>,_YQ_'X 
@4#(AAV_</$KZTIWU J<BLZFM.]R1#LI+Y'(BS)K@X%H 
@8*)SA9V K*UVY;8&Z;FN?X/ZX5IQ>:2P1SNR;%-^4"8 
@G8Z7%+&W#7&W;ZQ0+AMP0*L>/I5_)Y=SU;>_0\2:X$< 
@N\K2[A]2I"&B-#QLW,_-?>6QOX^_6_PTF_@P#[Q39]4 
@XZE+X&9>U&B0[=3!=W"G[8Y,U!K;!/4FS><$4365<,D 
@:VK2F4]MV((3WTQD/33W*IM2T?OS_JTAN2XZHY28)W( 
@ID7[@HQO+3'*T?QP$9CK.AALNW4>6]D^'/X.K'0),Y  
@YU#MJU3-98D476H6PVNFEH*_@<7*$7BD+RELTET!%B, 
@'] O M\UH'2L:],H\4!H/==!MM:J$<YWPY:1"Z42']$ 
@CE3"<DU";N?/(MQW:O^6[>J3@Q6P)(1 1&>\9]?X,S0 
@6G:9 W\E"G1_Q"7+O'I@)'.UW8Q(!5]<ZSM[IK^LV<L 
@A6& LF+<_OVQ7.1R$V/W6EFC9JD/F.]Y_K/1]8/@#.$ 
@&^+8TZ4N@XFT=4,J]!<3HZ%8-:$#ZC\EXJ 8!+:H3R  
@%M&OJMNP+GXOF)81_^'463,UD<:GZD.** HUR+/"X.( 
@P0[Z!^OKX;("&(9;Z!.KCGX?7RW<NMM#G,OTK5.XK38 
@*[\>XOW]!5 8 %1!GZ*50^2N(4I*Q'UHIO+NT4'&*(L 
@_\P$2/V=@?_Y)*#+XK$PS_F4)U7Y<8&/GPP%^W/L<#( 
@6ASNG0.K",]1/X;1NDI&J!]J3Y(]59X[;/A]IAD#FD$ 
@##4 LW@S?RD[['.$VB)$?N-^_^724TD/SNCEEU<'G#L 
@]Y U'S'F\MD,C("PY8C34/0+^WLH/]2G>X_46=>JB&< 
@F%!M-IRL/,N'R.+(V,*"6Y'YXYL^GQ?#&Y\.1]>][3< 
@HM,#E\*M@GS6;K,7,%6?(A&H@7)WYPAR8\K%,0HKXRP 
@+_%C?]G]ES0BQ0PP[RD;U,2"A*[,O,DPK.%<J9$:L:( 
@$5^124:C;O3&/I_9O=H$OLEU@),6T:V#H$(-!93U;P@ 
@FB,4\:4,=&]?%O1'*$>#= >J=_2;W)4BH-F)!<R",Z8 
@;V:<L:"S\NDWP0@-Y!WU.S4^\_,U%R?FCT!,50U)R)8 
@B4&QO[VX0^(&8J$,OHO!"BQI6Q53RGS+"!(NC3OJUZD 
@"Q"Z8D;'^H -7<T'2%1+0 X<V IKDZJ5#[]L1?WJ.'$ 
@NW#LZR;@<F0]9U )#E##W,Z8LC+447!Q1A9RR!R,7M  
@UY%["PDV\GCYK(9->MD:G.3; Q@!H$^C^I6 8'40/8$ 
@H@DVVT-C82=-#[G#5>*GS8JFF8ZZ=9P?=<[H7-H,7O0 
@^APU8F@QSB4 /5O8&PNA0_T*)[7SN/(C[U$A/*VCLP0 
@\JJTW& =,4\."Q"2SA*!8-#=O#R4[8 N?B*F#S %"L$ 
@AOT6%D'G(RJ_OH*[B_%.W;T%AS*"/,[EM#K!NS61K(@ 
@[Y7J@"G,((YZ%8;354=:O=]<2:/_S5[>ASOV<,1)>W, 
@,BC#A!SV/(.3.D!*S*3 @W^*+E]I^4/Q3C@I9.^(D$< 
@,SH9FW7#I2XS+[ML7,+'<B9K:)I3Y =.T9D29^VX:UX 
@F4$_9_5S]FBJ08XP<O#-+ WO@]=)8PWY3APR$Q5,JKD 
@>],_+L;SD)XVDBKZ'A_!\9=_JI:5SX+[UP-G@?9*'14 
@O9\W^OK)_A_S8P/K0"O+-R;^*4NS2<=58?U7?;<T*$, 
@%#&!LOH') :,K.TV"PWQ'S>F@0B_*-TD."#DZ%D6:=T 
@[Q)S-UQP!<$0(J?1YW5:AM2POL-9##YY_UNV#2P;/FD 
@J^0GR.=DY$S<U30Q:Y-$<G_U["-KM7=]/^/V]N++!$P 
@"/1HK[FX[<5"F/VHCN-#KIN?EYAUX(<XA"V/Q,! 3)\ 
@RWT75I^.1V&52YTD*J\*&O61/B"@Y-QR:?TE-JOI1A4 
@J'=T>..B08&1'T C(7PY83Y*%"+'3M:88;1J8Z<F3F@ 
@*EPP#W&XQ3[>(2+?IX$/2E(UON,AX6^-7_>A@&:146  
@.P3]+LPN5WG!?80PM;CL2D$EN?R2=ZBBC3H/:9D]_&4 
@F!F)M/G/4&UK](!SY;$!@A4'[.CL.6C$5HS4RD?O_I$ 
@2;A_65,E>;5$R;QCLZ1:41U0H;HC_:IY?QLCL8-RO;  
@_W;(N;+M^3X.ME8J8 GJ<3^+Y.98@^H69!$CZESHY)4 
@1J>P4>\ZH"S"4?8R)@_.P=,?JX<L.LOU8$ '8]^X[>( 
@V1QN9OK4I4%U>K"0H9&^N9$$IQ8<E43O6X;9@G"'F:@ 
@M(:8+C:V->M2\T^/WW-R$D+&D&7HTWK,%%!:VR\)E7X 
@&.P#R>^'.X_I)N AC"?!F\(_H3(?5?K+_:1*2STJ^3  
@90[F#%?ZOX0G0I":+L+2S/9 &LLPFN4"LSF9T)H[WOP 
@AQ932E-*VF[QXX)'$[1HU'Z7+)4&M/<0E'YN_ZJT) 8 
@V)@">A[T)[SIF?*VSXM.5:$)SC\A#,)918EBK:,O,]< 
@LG=U^\$:%"BZH [:J-O!CD^]KX=A?,:3V$>_+H8J+F4 
@S981X-!>?L\KB7$S5W,O2_6A3R:I6!;>4$#ACR;+55( 
@3<4(UOB6[Y;B\]1(".(DQ(6ZX# U8-V YC1RU7@@$-( 
@#%-28%7@RI<PY%\K'FU0]X].-"ZP/GL.+> ZQ\[A]V@ 
@<ZQ#4W^N&"QXJK !.VYHW[@U;5?BKIU@]=9NJT[HH., 
@99/:T:0X)3K\[-T,*HU.R#UP,!(QCKQ2797O<CKNR7, 
@EK_']+%/7RM>MM8:AY-<[?1KI7:-+*]IM%AH%]>7=C0 
@MSQ71Z[FG!$]325RGZ2+)14=&_;TRP;]++HRP#3Q<*@ 
@S3\^'I;[W[%#"VX>]4+2$Q+G:31Y(GQ<T$-%Y]?DIW@ 
@+B6&-G>?DDYHS6#P6EDR',V_E[1P3>J^8U] X-5JG8< 
@.M.$HY\28'=QOR)?L'>.,F]%(/S.Q^W8RBN3X-;MEYL 
0SF&W=Q</2#KUHREP6?*0FP  
`pragma protect end_protected
