// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 03:42:19 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VrO4z4ZvhdoPuUyZhmFW6ThCKYFWTOg5kCA6VP7uIRd84doTMCXEIkhKrRDN9+N6
2X5kiKfjFDIDiedvY4kr2QpkC1jUOovCz19J+DnRpEGZlEVQRwC6u457tukS7xE1
/posNM9+5n19f9DtfS1jP10an4NMl/EC6ni/yHOLDTQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5184)
Fw+LTbl3Rf4Pvk2nnRXvi1P3jNm7vGTa30l7pvW2zTI6lmfbUm5HJI0ydobP6zwA
f8SqIoW05/L4N3adkhWKTDIVQuTLVDzSIQF1qcdeRz3s4JoYRFaurZ7GjtsO7rKk
P68KDQmwirqqqaIirfwQAJ6ylaA2vNYpnoykewLYoEyyvk8oH/A58SBBIsS+fWQn
Rzk2yJflpP+bvVN1vno5vTi3ckksezD2hLLMgq+jVGbHFWXsg2KXOC2113uc2WsA
1lDtocGJfaW7iu027wcdZrsjWGLqEbh5w41QCptZN/p9maAkHfCk7rcoXEj7QIY8
aBV9aDDiwII5hYQvzog7fMvAHehvseL0M9Gjmeth6gtce7OJwtNmPs3Xmwa4Kn25
VnjY+7h/iYZ60ouIihG2Qk+vBqEcLIBCqS/8sURXeOMyMYpfNft+wEacc1MkBVmu
tmWebJhTqAlvNw4FAudnB8vrr4NOn5Je8z5LsGXHI1yTMtRodIyNol7i0UHDg2zF
xLaUtKEQSuHd5VPu+LztrVEbjCRYB65wJtI7UD+K1H/nGF8ttHmvXS2p9H0BJjYO
5wSlOqLhPBl3nqgsNxx7U209LfArd/OdTcGBtosCf3Ruj1EoS3nHkMsq8VOnh40V
AXr7Ea7e1TMobYZn9aYW1xM7IflW7ockEnjdfLozin9kmI8E1uc7q535ZYakJ5C2
YjSGuMA+P+Gfv28HavvfzqedU6v3ABhXWONAuwW+DNTwEaBHj0lBZm4vVBi/e/nD
lcVn+KH02OkahnIBSEbzKIOYgo8UFFh9NZPEBZ3dru554BxZKEt8E71T8qUWYFX7
/veJG/gkcobZr3zthxJQgcD/N8tYOQHsdeHk/ucdlmf5+1YpJgTFldCrPkDEw1A2
oBNIHZzjlYvCZ0aRx+qwZEUHFDu5WWdIfxkZDaWJoB0bnm8SbIJRJSo9IkvacMrT
F4nX0zPEdKPMFiXpOxIvJ3zyxXH3HWTdysTCqN6wvuNz1XO3jJDgBqMIjl7ZVMPj
7awwvtBa9D1JZHT5clMnqfQF39ViFcUPn1Z9Ld+sMEK53mPjD39ih6W2cjBj9Pso
egqrKrbdGqDQltM+qb31J5LopI206rqUHfjOuaiLgwEp1qB6/qTDu4m3OjsS2xSP
4ZQkHh3Nca53GQb26KUbD3zOvaShP8rlKdL01umhmLIhyv1q3g6l86R1wzGxl8qL
GfLvpoVWWnxa0WkdaRctGnkdkom4VgGlpa0dsnLoAyevVZtBTGsUvdIB15CVvVqt
XsbGK9sqGWFQu/FKiQi1PK2JDEEXXTo6Oz+1ExQYgBrsRxeFG0Y8Ze6+KS98fRWG
fvzKp82xtBcVIwmfE1w3JdTVdGI2cCdHj517EoAocBZP9mK9QKS32cyWYdC2/22O
EkWVPGawMe0WT8HkJk3ITDClDV9kXOkzY813J/omII0nIWdDJ/03++Bl06I0X9jv
xcdcNWSRHUywzh2WQtZGIBLzLxAWhwelxQINy9/ZZIDXDSbABzfVd+esa3vWqxcm
HqfeiyqpXUs5QGkHLqtddK2y2AY4pl7xdfVa9Th5GcHgkuU7FWXb+dgbFbTTD23Q
/dxaxlfzodxlVtagV+8E+1qVLMSVDNdN5J3ezLrrbrerbrKyXYJsWCFg6OM7pPYg
Pv5sonJKX+OsFWCMiTuToVvNGPCuANGHBYCkSS5toSIxLIStaSJYjMT6PVRVcy0k
38cglvqjS2UIdLl57xoVR96G+Lk5KTeTtOVJHAVYaS+VwqDAzTsn4g6eCfqX4n1x
tMnIUmuvFqn1s0EZ1zIbcyGTTwH6sw2/EEsD+dmubAls+bk1T7tHaN9pHZVoRoZT
E2fWhU6+zZLNZQkDJAVHZux36Izoxb0IN4MI+6NfaNDXQuPGYgHog5KCYWXavi46
WFnCgHEI8GhdT8XAYxM1m6nf/+j4bNDAdhC9SRWTJ3qQ9fyg3HZ50rrW/faA+P97
gam1YZJYQYSUdamLKNUDe1mdpH4aNrWXksVdcwhKrFAaR5Z2d89a6+Zl6DyL1RBy
cwQyyp3tF9DDQRxr+UiTYCgRIhYOrXsY2bJaYXypr6EwgCxWQQwu1vZYiZ6vYznr
dyWNhQBB7zOfiZzKJwkib1AchDch4j7E9Mgy408tFrWtDkJzV5WTET7Ihtocrt94
umCgbXD58o/8vPnPSsylxhq01RMCaRZt7LqZDMuARUR3vKe8ppl1tCEKdyMtHwJ6
3eL3trrY/zET4zMR4itN1MsC0WISP+fLJN9eVLDF52I1LnWYtlzPQR2zkuY7ZhsO
xx/yx1ibAuyZFKJoVbfiyW5tIHhKhstpew5lLgX2rkPfAaxUj10e+tU2vkOtGnUs
GnbdWRIfSrlsB89rqpKj/SqbvTCE01PClH1ctACA4BfTlKdOUjlGKOb8V91lFLYz
dZGcjko1Q6xZe5YSeBjlxGN1im3A7ImIrQCZj9m/KQJZLNl+M4t+9KbxzlCrZkhg
NlbjCRls0lsqtGeqXPURWUmJ4ac89nTjNLp4O8iPZAdy3MykNMD5IIqEwOirgaqz
5rq+gCP5l9XzfVvzclATeEgI1rN/F8mOPz+99iIIw0zjHZR/4MrALupoAv45OxiZ
mEjE8zJg43EyFGSsopritM/eWnuwQTFSkZE85hC/RCpAKaplKepMC/iH9XLzwSTD
RHbnVvok1oslgmMa40jKPcJfD2OFBX6g9fgNvBdUgKWw3PjqLPqgJYAj9qAQLAv1
gLHpSIPUvo/PJW1CLEsQHkNeuUYlC5WgHXAxWep64qUgj43WTh6+DZYSr7BBTzTD
U5e/FxJU/xIgPfXaeSKks0IVijPvwrvVYJeGTRp0gZglVt8Cu/bmTPN4krwlrhmx
f8Di4Qx9OodP9M6qgHvdOgCWO8zsSbe9kMnzdU14fx2IsdC7euFqstwXkrg9If9+
3PStolPIPeiJCw8GPUhxDGIVXlGD30xncx3t4a/CoGwaoPJ6yyk1lruC4MwmzM/D
2KDVXw7IEaKjrLya3qneBSfYEH0R290HbovWI64FKZt8jGuZzIh2cs2N6I2fYcOF
6N0YftHC20mfk1fpytsq36ZXedq0snpUGc9AR7tHY/2sCfOj8pukh+E353Gg6VMA
Ug7IB/yNsL+P3speOOD0BJ756MvpdlJ3yWO1LXV9kiiZup1jtLwdZCdFK9cvy31A
kJA9CWEwoTIbpvB3zQPkmbRud6VvynlWHgwVl6AWnaBtSroPGUriLSfUpqS4QTDJ
rWktUecRShQP1dC9idbJuJMhol9KIAQWXRDtMuog4mmak7sie10xNa9LR0PVqbuc
ZXLDhzkGac4lpQ7XgJBRweFv0wJJ2+JptP6+Bq0+yxkybJwdlfXkJUUijPuBVzVI
X7yWNnRAivSlFvDDWQPaDvtHJAaEGEUgrer1bmE9wnZvyv1UvDm3YEhQcHHU0LEZ
J5jcDG2+jHKhS98YSfXHR8dmSX2XlhyY0NNrmp3CvfhtnTUglxsjaqWd55jB4Irs
XozKPwEu78zsDWGJK6AR34cuwuAr8BPrTlDY9Zn6tjwsbD0/Qb2BLZ6BTPYINn/n
feFYIfxQfnIyk3KhtKGDN3XgW0niz3AXjwQQ0UspH4x7WBY7JU0b1eWuFazEkzzY
P6fTeeDECakn2jxSUiaSVc6/YpVAE2aV5AjLgdNW68qYRxuQPCOrgY+Vb4WgLeav
1TIXM3VkOplke2gFF9Ly2hxLaTPkZinDef/BTLYL8bEYx//cerYo10Vtxnw9hE1x
jWRhfhlG71vwZYRfFyqlg2QQAsIZ5QzhZLN9w91T+3uHhGRvYLsTjNz1idGW/6SO
dFxogr2WfRTPM2dmbvjUDw8TPhT4gY+lgyau06y4SvzbNO2rKCvW3gmksKSryu4f
FWXCtP/7ZwPNwP34CkVOrYU40Cq4Gvf2hymxAot5FrZ1yTeXTUJHQ1WCCHwnFZBS
41ljObxU/ZzoIBESfS01v4fsKwfRP73IC8z5Byj79+Rv0PEEbWJSrDPIpTC7/Vlb
5Y8ZqlLewDzQtN1YikLKkBBmbhHtvgEzU942OtBHNGI5cece81j2w8ONrduesjEL
K3T7iS2Q0koO0zinF352WyyUBclMLBriMVlVHeR4N0kI/QS+SiWRnxekSCW6GjK4
LpM+fAMM2rtyayOOTXIz/K24qkZPUCMag3KAQxYNHxgFk5amKRsZJdwznTyahHK+
svm4vksBg0LONqWXNYGO9I5h3WhO2cn0qiGK/AuAYuUwMgpDyXyG4DQskVN3ca6K
XuuKhGJFy1Gwx1nAOFdanH8H8BGTf2MZDvy55E59Q1tmKCDqmfwdxRGLtgEhZ/lO
QRMYqkZiiMNd1i6OBBt3qQrtcI6Qm8loLE7YtOlruxBhrDFdZA/1+dsbhRAaI2cF
7HyYKJrvM4B9sGFennscSO+6VGP6lMzCa4qpZPaFiF3nMFXPSNDvKemCvMVyu8SH
PEd1c3kaXkpITA3odwG/rqcASXtREnh+cbAxvZnCLRpcmBRPa3lPeWlSn8wJZIaL
sygDw9SU4qkGv8wqSiTGsm8DIBdiJjB1cLikjO2TuBCh8Wbc8OGhx92UGR+Vl7lL
vEm4f6Tw5ZXfXRmP9QOcvyXTbmmw7uG4qYct2/V2fQScUvrwCd8TnVGDlq5Dj4ge
ET0xcw2WKv+wiNebFptBlge8EIsJ702eyiSLAlQN0W9r+2+1GVLfIutnpvDJ7t1w
Aj8DjJvbRfDZZDB5dyVqffQPgQfOtoOpHzSKO23cGJqOyWUse0sbHYMtpUpCLstt
xFrsJU0wB1dYsZMj+Qo7+K7yD61+P5gLQqtfl1sFiReiMskK/3FZ1FSlDp/dnqkS
nQDclchBqxvR+zX/q+670iZGlVf8kALoXatT39VEBYg5MbIHJUP8igzIyd5dHGLi
AvGkocxv5+RCM4+coHOlFF06wC7NH+CSCrf4g9kRPZ8tiRzj6SViyM6Pjqxcvodz
595j4HoZW8DeBzXn/AjyKM/ubSW/hxiQM2r9BYW8A2nUGDxY6DfGtBkN0c+xRqQA
vHWquby2ZEwNvCGFAJt4WV8l8aPnABE3OyzH9WErhNrWBAlLC071F2R5/5DfA6wB
z4CQfWVe8gt2gJrvBSWQoYFrNaOPQDtaQPHgPhyATD+TqTTfPanfa7C/zHziJtwL
7QZYuOVotRFqzoFbvzg2p+ctSt2gnU622kLsO41IsKIEhxk0Ydw79pkKRV03QGdt
gA0eKyHpz/ADKvXrjV6x4kcYCZ7h3vjI3mKiLiwqX26rrdXcrIgGMxR+0IwUCDVr
a1DioYlAGa+gx2U2EsfzDjbfw0du8jNGa9HllAMADtCuEY+HDaM4gnX/WXeD4H8B
NuURFzyCqmeg3HUtmRh2jfV0EmX2VgIe0o028NdH1bEbln7+EPtn/SHgLaXjyXAg
leeG2XXcbhVLnO7D5P7FCBtRUtpngnnIlm+YcvaoHYe52bPeSoq/OpByTXMCZY/8
Lf/A4hiQN7kbhnFZYIRNr9TjGFzlafi75TW10g1v9A+u63nFMIwjrUz86+RH2xkU
dDVVXum261g+cgObAhl0T5akw47LXEYtcNDYf+0jiD6L7pp6r2jymvAi4o9PtKC2
mw09vOzJ2DN3uyuDSnOZ4tGKVc1/5wAMh/pS4AncA8NQ7iFv4+FG/S3yjuTLfhtW
c0ULpuEh7W6w0C5j5td8QevtKfu+arvkEg9FPxrc0rCBKkm02aN3MsMjsmKED9Sq
o7pqR6MC6huP3k6JBNipIZ57Hn0ezKw8EpXMMAiJQQy5nRwh9OK02upMKMJGZ1So
p3BdAMTWaAK0W1sIicUtO15jXiKMV6Al24k19Lcey93p5gzvJuPM1DYOTW/djfyS
I8nrRB54e/6OSaH0h7Jip1ked8k1xvs1IeARXlXok0hxNKYMOq1gAAQMCGOgGzrH
Mw4U/8edmxQgqj9bh5MsgeH5qBCSpjV5HobKvHeQ6+rALhvr7Dyx9BiDF8sXQbQR
79U3/db2zn2Izh0TWolpNHjLQ0HPKky9b6QLZnHcAMiWH4J5A4jcgp5gDi//m4IT
NNl5UsH5d3nWTtTkCfWHs019HzOi8nFOF/sXquLjc4I4aGKFjv03ALT5udVlmySQ
zDmW2n77Zs9KMIkMqRNBWEDQ8wgZ7JN1QfCKdOyCfemKkj+ftMjbL6H+jD35iydY
SG9sB+/qPgsy6GT7vLlOfRxPDjAWBCyFftaE89R9DmGKZQKDsOJiq6CXEnR7OvEh
wzkoiB9OqhEeDpeujC5JR8Y9DEWrZXc0d0OYqsTFjDyJsPeN/sJYsmsmGbVxN7yQ
SUctmRGVTh+vrHKWF9zb38Ed7QgrkNokxRsHbGX3+1hpmrH82cuPjT4DqwkQ+wp4
BN6LarKa7maxBSGCO9MC0FjTDgq/2UBqM9pq1zXRUpZSaTrVswUuL+ULuulsIWqI
4DJkISRbpxZaeupA7xoUfLh2a9us9kAvFRzV2Nav15qCxRlYk72ODidT8xH3+mJ/
gJkrHn3fA8k7jtle4zNobgQR3VZL+hDapfaSotYfmC+5CaQRucKFXyOlghhjqfwS
3dQkcqDjt2j8Krw/S+W4n6n92vFZ2JWr+Z0in+DSgav8UyuujTW6U5xsq8hLk2pi
6XhiEvwb3ixNrTZIIiYBlDPpY0ohNvYKMGmwnMSUf5k7CW0PbYBQ0DIE0h6PaAUw
ZwOehmlBSzgpNma9efX1cH44a1qUG8sKGw/3oNxmutawPEtwkUIdmAsgpv+AeWMQ
V5X7b2NfrCcqn4rpD/k6MWU2KudFNxOSGce/BglWr80Kom+VTdqtXfRMm72zcjbo
gQ07dUKmGFo+4TfBfgqnGsdUM9NTXRbbfkjmHNYFj+ChXHkOBgnUY2Ywv/+nBNQp
`pragma protect end_protected
